/*******************************************************************************
  Copyright 2019 Andreas Brokalakis
  School of Electrical and Computer Engineering 
  Technical University of Crete

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.

  ACKNOWLEDGEMENTS
  
  1. Some parts/ideas for the code written below were taken from the source code
  provided by Supranational here: https://github.com/supranational/vdf-fpga
  2. This code has been written as part of my submission for the FPGA Contest 
  organized by VDFalliance: https://www.vdfalliance.org/contest 

*******************************************************************************/

/*
	INITIAL CONCEPT
   -------------------------
   The following were the initial idea behind the multiply that was provided by
   vdf alliance.
   
   Multiply two arrays element by element
   The products are split into low (L) and high (H) values
   The products in each column are summed using compressor trees
   Leave results in carry/sum format

   Example A*B 4x4 element multiply results in 8 carry/sum values 

                                           |----------------------------------|
                                           |   B3   |   B2   |   B1   |   B0  |
                                           |----------------------------------|
                                           |----------------------------------|
                                     x     |   A3   |   A2   |   A1   |   A0  |
                                           |----------------------------------|
      -------------------------------------------------------------------------

       Col
   Row     7        6        5        4        3        2        1        0
    0                                       A00B03L  A00B02L  A00B01L  A00B00L 
    1                              A00B03H  A00B02H  A00B01H  A00B00H          
    2                              A01B03L  A01B02L  A01B01L  A01B00L          
    3                     A01B03H  A01B02H  A01B01H  A01B00H                   
    4                     A02B03L  A02B02L  A02B01L  A02B00L                   
    5            A02B03H  A02B02H  A02B01H  A02B00H                            
    6            A03B03L  A03B02L  A03B01L  A03B00L                            
    7 + A03B03H  A03B02H  A03B01H  A03B00H
      -------------------------------------------------------------------------
         C7,S7    C6,S6    C5,S5    C4,S4    C3,S3    C2,S2    C1,S1    C0,S0
         
      
      IMPROVED VERSION
  ----------------------------
  
  Since we actually want to do a squaring therefore it is AxA rather than AxB
  then we can make a lot of improvements.
  
  1.
  Basic observation: since A and B are the same, in the picture above notice that
  for example A01B00 will be the same as B01A00. Therefore we can seriously reduce
  all multipliers required from n^2 to (n^2+n)/2
  
  2. 
  Based on the previous observation, in each column the terms, for example,
  A00B01L and A01B00L are the same. As a result, we can shorten significantly the depth 
  of the CSA tree, by using only the upper half of the grid and using all numbers multiplied
  by 2 (which is not a true multiplication but a shift), except for the numbers in the main
  diagonal which are unique.
  The result is that in the tree now we have to add at most n numbers instead of 2n-1
  
  3.
  Reducing the tree depth by as much, means that we can follow a much wider multiply strategy
  without sacrificing clock frequency as the critical path becomes significantly smaller.
  
  4.
  Problem: the above work only for squaring and NOT for general multiplications. This means
  that the strategy described cannot be generally applied in the reference source code provided by 
  vdfalliance. 
  Solution: It is now possible to complete the whole squaring operation (for all elements + 
  redundant elemements, i.e. no segmentation) in 2 cycles and the synthesis/implementation
  prove that this can be done safely @250MHz. 
  
  Note: the drawback is that significantly more DSPs are now required.        
  
  5. 
  The code here unifies the next step - i.e. the CPA addition - using adders in DSPs. The result
  is available in 3 cycles (Cycle 0 : core multiplications, Cycle 1: adder tree, Cycle 2: Carry 
  Propagate addition).
  
  
  NOTE:
  A custom C program has been written to autogenerate the code for the multiplier instantiations.
  NOTE 2:
  The code reuses the provided compressor_tree_3_to_2 with no modifications required.
  
  
  
*/

module multiply
   #(
   	//MODULE PARAMETERS
   	
     parameter int NUM_ELEMENTS    = 66,
     parameter int BIT_LEN         = 17,
     parameter int WORD_LEN        = 16,

     parameter int MUL_OUT_BIT_LEN  = 2*BIT_LEN,
     parameter int COL_BIT_LEN      = MUL_OUT_BIT_LEN - WORD_LEN,

     // Extra bits needed for accumulation depends on bit width
     // If one operand is larger than the other, then only need enough extra
     //  bits based on number of larger operands.
     parameter int EXTRA_TREE_BITS  = (COL_BIT_LEN > WORD_LEN) ?
                                       $clog2(NUM_ELEMENTS)    :
                                       $clog2(NUM_ELEMENTS*2),
     parameter int OUT_BIT_LEN      = COL_BIT_LEN + EXTRA_TREE_BITS
    
     
     //END MODULE PARAMETERS
    )
   (
   	//MODULE INPUTS
	input  logic 			clk,
	input  logic [BIT_LEN-1:0]	A[NUM_ELEMENTS],
	input  logic [BIT_LEN-1:0]	B[NUM_ELEMENTS],
   	//END MODULE INPUTS
   	//MODULE OUTPUTS   

	output logic [BIT_LEN-1:0]		reduced_output[NUM_ELEMENTS*2]
	
	//END MODULE OUTPUTS
   );
   
   //some local parameters
   localparam int GRID_PAD_SHORT   = EXTRA_TREE_BITS;
   localparam int GRID_PAD_LONG    = (COL_BIT_LEN - WORD_LEN) + EXTRA_TREE_BITS;
   
   
   //DONT FORGET TO ADD SIGNALS REQUIRED HERE!!!!
   
   //please check comments below why this formula is used
	logic [MUL_OUT_BIT_LEN-1:0]	mul_result[((NUM_ELEMENTS*NUM_ELEMENTS)+NUM_ELEMENTS)/2]; 
	logic [OUT_BIT_LEN-1:0]     	grid[NUM_ELEMENTS*2][NUM_ELEMENTS*2];

	logic [OUT_BIT_LEN-1:0]	Cout[NUM_ELEMENTS*2];
	logic [OUT_BIT_LEN-1:0]	S[NUM_ELEMENTS*2];

	logic [OUT_BIT_LEN:0] 		grid_sum[NUM_ELEMENTS*2];
	logic [BIT_LEN-1:0]		reduced_grid_sum[NUM_ELEMENTS*2];
   
   //SIGNALS!!!!
 
 
//CYCLE 0 

// Feed the core multipliers with input data
   
   //First produce all products
   //Instantiate all multipliers (each multiplier is a DSP48E2 but from the slice
   // we only use the multiplier and not other functionality. Remember that the 
   // product is registered, therefore results will be available in the next cycle.)
   //Important: since we are basically squaring (A = B, dont care that both inputs are set
   //independently, this is for compatibility reasons), we dont need to compute all different
   //products (the product for example A1 * A0 is the same with A0 * A1) and therefore
   //we need instead of n^2 only (n^2 + n)/2 multipliers, where n = NUM_ELEMENTS.
   
   //no easy way to autogenerate the instantiated blocks :(
//A0A0
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B0(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[0][BIT_LEN-1:0]),
			.P(mul_result[0])
		);
//A0A1
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B1(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[1][BIT_LEN-1:0]),
			.P(mul_result[1])
		);
//A0A2
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B2(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[2][BIT_LEN-1:0]),
			.P(mul_result[2])
		);
//A0A3
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B3(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[3][BIT_LEN-1:0]),
			.P(mul_result[3])
		);
//A0A4
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B4(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[4][BIT_LEN-1:0]),
			.P(mul_result[4])
		);
//A0A5
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B5(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[5][BIT_LEN-1:0]),
			.P(mul_result[5])
		);
//A0A6
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B6(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[6][BIT_LEN-1:0]),
			.P(mul_result[6])
		);
//A0A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B7(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[7])
		);
//A0A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B8(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[8])
		);
//A0A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B9(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[9])
		);
//A0A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B10(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[10])
		);
//A0A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B11(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[11])
		);
//A0A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B12(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[12])
		);
//A0A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B13(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[13])
		);
//A0A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B14(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[14])
		);
//A0A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B15(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[15])
		);
//A0A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B16(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[16])
		);
//A0A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B17(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[17])
		);
//A0A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B18(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[18])
		);
//A0A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B19(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[19])
		);
//A0A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B20(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[20])
		);
//A0A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B21(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[21])
		);
//A0A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B22(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[22])
		);
//A0A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B23(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[23])
		);
//A0A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B24(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[24])
		);
//A0A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B25(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[25])
		);
//A0A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B26(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[26])
		);
//A0A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B27(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[27])
		);
//A0A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B28(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[28])
		);
//A0A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B29(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[29])
		);
//A0A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B30(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[30])
		);
//A0A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B31(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[31])
		);
//A0A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B32(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[32])
		);
//A0A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B33(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[33])
		);
//A0A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B34(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[34])
		);
//A0A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B35(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[35])
		);
//A0A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B36(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[36])
		);
//A0A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B37(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[37])
		);
//A0A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B38(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[38])
		);
//A0A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B39(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[39])
		);
//A0A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B40(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[40])
		);
//A0A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B41(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[41])
		);
//A0A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B42(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[42])
		);
//A0A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B43(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[43])
		);
//A0A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B44(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[44])
		);
//A0A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B45(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[45])
		);
//A0A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B46(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[46])
		);
//A0A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B47(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[47])
		);
//A0A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B48(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[48])
		);
//A0A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B49(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[49])
		);
//A0A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B50(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[50])
		);
//A0A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B51(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[51])
		);
//A0A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B52(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[52])
		);
//A0A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B53(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[53])
		);
//A0A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B54(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[54])
		);
//A0A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B55(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[55])
		);
//A0A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B56(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[56])
		);
//A0A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B57(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[57])
		);
//A0A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B58(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[58])
		);
//A0A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B59(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[59])
		);
//A0A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B60(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[60])
		);
//A0A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B61(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[61])
		);
//A0A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B62(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[62])
		);
//A0A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B63(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[63])
		);
//A0A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B64(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[64])
		);
//A0A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A0B65(
		.clk(clk),
			.A(A[0][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[65])
		);
//A1A1
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B1(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[1][BIT_LEN-1:0]),
			.P(mul_result[66])
		);
//A1A2
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B2(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[2][BIT_LEN-1:0]),
			.P(mul_result[67])
		);
//A1A3
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B3(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[3][BIT_LEN-1:0]),
			.P(mul_result[68])
		);
//A1A4
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B4(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[4][BIT_LEN-1:0]),
			.P(mul_result[69])
		);
//A1A5
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B5(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[5][BIT_LEN-1:0]),
			.P(mul_result[70])
		);
//A1A6
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B6(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[6][BIT_LEN-1:0]),
			.P(mul_result[71])
		);
//A1A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B7(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[72])
		);
//A1A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B8(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[73])
		);
//A1A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B9(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[74])
		);
//A1A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B10(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[75])
		);
//A1A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B11(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[76])
		);
//A1A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B12(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[77])
		);
//A1A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B13(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[78])
		);
//A1A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B14(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[79])
		);
//A1A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B15(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[80])
		);
//A1A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B16(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[81])
		);
//A1A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B17(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[82])
		);
//A1A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B18(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[83])
		);
//A1A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B19(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[84])
		);
//A1A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B20(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[85])
		);
//A1A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B21(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[86])
		);
//A1A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B22(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[87])
		);
//A1A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B23(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[88])
		);
//A1A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B24(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[89])
		);
//A1A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B25(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[90])
		);
//A1A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B26(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[91])
		);
//A1A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B27(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[92])
		);
//A1A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B28(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[93])
		);
//A1A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B29(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[94])
		);
//A1A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B30(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[95])
		);
//A1A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B31(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[96])
		);
//A1A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B32(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[97])
		);
//A1A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B33(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[98])
		);
//A1A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B34(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[99])
		);
//A1A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B35(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[100])
		);
//A1A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B36(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[101])
		);
//A1A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B37(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[102])
		);
//A1A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B38(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[103])
		);
//A1A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B39(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[104])
		);
//A1A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B40(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[105])
		);
//A1A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B41(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[106])
		);
//A1A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B42(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[107])
		);
//A1A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B43(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[108])
		);
//A1A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B44(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[109])
		);
//A1A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B45(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[110])
		);
//A1A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B46(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[111])
		);
//A1A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B47(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[112])
		);
//A1A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B48(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[113])
		);
//A1A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B49(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[114])
		);
//A1A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B50(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[115])
		);
//A1A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B51(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[116])
		);
//A1A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B52(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[117])
		);
//A1A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B53(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[118])
		);
//A1A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B54(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[119])
		);
//A1A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B55(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[120])
		);
//A1A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B56(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[121])
		);
//A1A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B57(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[122])
		);
//A1A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B58(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[123])
		);
//A1A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B59(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[124])
		);
//A1A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B60(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[125])
		);
//A1A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B61(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[126])
		);
//A1A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B62(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[127])
		);
//A1A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B63(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[128])
		);
//A1A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B64(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[129])
		);
//A1A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A1B65(
		.clk(clk),
			.A(A[1][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[130])
		);
//A2A2
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B2(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[2][BIT_LEN-1:0]),
			.P(mul_result[131])
		);
//A2A3
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B3(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[3][BIT_LEN-1:0]),
			.P(mul_result[132])
		);
//A2A4
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B4(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[4][BIT_LEN-1:0]),
			.P(mul_result[133])
		);
//A2A5
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B5(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[5][BIT_LEN-1:0]),
			.P(mul_result[134])
		);
//A2A6
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B6(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[6][BIT_LEN-1:0]),
			.P(mul_result[135])
		);
//A2A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B7(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[136])
		);
//A2A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B8(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[137])
		);
//A2A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B9(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[138])
		);
//A2A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B10(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[139])
		);
//A2A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B11(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[140])
		);
//A2A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B12(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[141])
		);
//A2A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B13(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[142])
		);
//A2A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B14(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[143])
		);
//A2A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B15(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[144])
		);
//A2A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B16(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[145])
		);
//A2A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B17(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[146])
		);
//A2A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B18(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[147])
		);
//A2A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B19(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[148])
		);
//A2A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B20(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[149])
		);
//A2A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B21(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[150])
		);
//A2A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B22(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[151])
		);
//A2A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B23(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[152])
		);
//A2A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B24(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[153])
		);
//A2A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B25(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[154])
		);
//A2A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B26(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[155])
		);
//A2A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B27(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[156])
		);
//A2A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B28(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[157])
		);
//A2A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B29(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[158])
		);
//A2A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B30(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[159])
		);
//A2A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B31(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[160])
		);
//A2A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B32(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[161])
		);
//A2A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B33(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[162])
		);
//A2A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B34(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[163])
		);
//A2A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B35(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[164])
		);
//A2A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B36(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[165])
		);
//A2A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B37(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[166])
		);
//A2A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B38(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[167])
		);
//A2A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B39(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[168])
		);
//A2A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B40(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[169])
		);
//A2A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B41(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[170])
		);
//A2A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B42(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[171])
		);
//A2A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B43(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[172])
		);
//A2A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B44(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[173])
		);
//A2A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B45(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[174])
		);
//A2A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B46(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[175])
		);
//A2A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B47(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[176])
		);
//A2A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B48(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[177])
		);
//A2A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B49(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[178])
		);
//A2A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B50(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[179])
		);
//A2A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B51(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[180])
		);
//A2A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B52(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[181])
		);
//A2A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B53(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[182])
		);
//A2A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B54(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[183])
		);
//A2A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B55(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[184])
		);
//A2A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B56(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[185])
		);
//A2A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B57(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[186])
		);
//A2A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B58(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[187])
		);
//A2A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B59(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[188])
		);
//A2A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B60(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[189])
		);
//A2A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B61(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[190])
		);
//A2A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B62(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[191])
		);
//A2A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B63(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[192])
		);
//A2A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B64(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[193])
		);
//A2A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A2B65(
		.clk(clk),
			.A(A[2][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[194])
		);
//A3A3
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B3(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[3][BIT_LEN-1:0]),
			.P(mul_result[195])
		);
//A3A4
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B4(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[4][BIT_LEN-1:0]),
			.P(mul_result[196])
		);
//A3A5
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B5(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[5][BIT_LEN-1:0]),
			.P(mul_result[197])
		);
//A3A6
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B6(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[6][BIT_LEN-1:0]),
			.P(mul_result[198])
		);
//A3A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B7(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[199])
		);
//A3A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B8(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[200])
		);
//A3A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B9(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[201])
		);
//A3A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B10(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[202])
		);
//A3A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B11(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[203])
		);
//A3A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B12(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[204])
		);
//A3A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B13(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[205])
		);
//A3A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B14(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[206])
		);
//A3A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B15(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[207])
		);
//A3A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B16(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[208])
		);
//A3A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B17(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[209])
		);
//A3A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B18(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[210])
		);
//A3A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B19(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[211])
		);
//A3A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B20(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[212])
		);
//A3A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B21(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[213])
		);
//A3A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B22(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[214])
		);
//A3A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B23(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[215])
		);
//A3A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B24(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[216])
		);
//A3A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B25(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[217])
		);
//A3A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B26(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[218])
		);
//A3A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B27(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[219])
		);
//A3A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B28(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[220])
		);
//A3A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B29(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[221])
		);
//A3A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B30(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[222])
		);
//A3A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B31(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[223])
		);
//A3A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B32(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[224])
		);
//A3A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B33(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[225])
		);
//A3A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B34(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[226])
		);
//A3A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B35(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[227])
		);
//A3A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B36(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[228])
		);
//A3A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B37(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[229])
		);
//A3A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B38(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[230])
		);
//A3A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B39(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[231])
		);
//A3A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B40(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[232])
		);
//A3A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B41(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[233])
		);
//A3A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B42(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[234])
		);
//A3A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B43(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[235])
		);
//A3A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B44(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[236])
		);
//A3A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B45(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[237])
		);
//A3A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B46(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[238])
		);
//A3A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B47(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[239])
		);
//A3A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B48(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[240])
		);
//A3A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B49(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[241])
		);
//A3A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B50(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[242])
		);
//A3A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B51(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[243])
		);
//A3A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B52(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[244])
		);
//A3A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B53(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[245])
		);
//A3A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B54(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[246])
		);
//A3A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B55(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[247])
		);
//A3A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B56(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[248])
		);
//A3A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B57(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[249])
		);
//A3A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B58(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[250])
		);
//A3A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B59(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[251])
		);
//A3A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B60(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[252])
		);
//A3A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B61(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[253])
		);
//A3A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B62(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[254])
		);
//A3A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B63(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[255])
		);
//A3A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B64(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[256])
		);
//A3A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A3B65(
		.clk(clk),
			.A(A[3][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[257])
		);
//A4A4
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B4(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[4][BIT_LEN-1:0]),
			.P(mul_result[258])
		);
//A4A5
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B5(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[5][BIT_LEN-1:0]),
			.P(mul_result[259])
		);
//A4A6
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B6(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[6][BIT_LEN-1:0]),
			.P(mul_result[260])
		);
//A4A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B7(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[261])
		);
//A4A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B8(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[262])
		);
//A4A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B9(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[263])
		);
//A4A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B10(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[264])
		);
//A4A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B11(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[265])
		);
//A4A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B12(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[266])
		);
//A4A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B13(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[267])
		);
//A4A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B14(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[268])
		);
//A4A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B15(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[269])
		);
//A4A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B16(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[270])
		);
//A4A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B17(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[271])
		);
//A4A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B18(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[272])
		);
//A4A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B19(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[273])
		);
//A4A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B20(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[274])
		);
//A4A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B21(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[275])
		);
//A4A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B22(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[276])
		);
//A4A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B23(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[277])
		);
//A4A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B24(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[278])
		);
//A4A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B25(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[279])
		);
//A4A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B26(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[280])
		);
//A4A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B27(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[281])
		);
//A4A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B28(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[282])
		);
//A4A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B29(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[283])
		);
//A4A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B30(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[284])
		);
//A4A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B31(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[285])
		);
//A4A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B32(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[286])
		);
//A4A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B33(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[287])
		);
//A4A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B34(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[288])
		);
//A4A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B35(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[289])
		);
//A4A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B36(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[290])
		);
//A4A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B37(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[291])
		);
//A4A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B38(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[292])
		);
//A4A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B39(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[293])
		);
//A4A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B40(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[294])
		);
//A4A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B41(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[295])
		);
//A4A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B42(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[296])
		);
//A4A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B43(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[297])
		);
//A4A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B44(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[298])
		);
//A4A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B45(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[299])
		);
//A4A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B46(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[300])
		);
//A4A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B47(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[301])
		);
//A4A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B48(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[302])
		);
//A4A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B49(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[303])
		);
//A4A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B50(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[304])
		);
//A4A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B51(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[305])
		);
//A4A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B52(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[306])
		);
//A4A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B53(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[307])
		);
//A4A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B54(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[308])
		);
//A4A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B55(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[309])
		);
//A4A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B56(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[310])
		);
//A4A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B57(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[311])
		);
//A4A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B58(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[312])
		);
//A4A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B59(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[313])
		);
//A4A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B60(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[314])
		);
//A4A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B61(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[315])
		);
//A4A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B62(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[316])
		);
//A4A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B63(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[317])
		);
//A4A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B64(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[318])
		);
//A4A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A4B65(
		.clk(clk),
			.A(A[4][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[319])
		);
//A5A5
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B5(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[5][BIT_LEN-1:0]),
			.P(mul_result[320])
		);
//A5A6
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B6(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[6][BIT_LEN-1:0]),
			.P(mul_result[321])
		);
//A5A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B7(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[322])
		);
//A5A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B8(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[323])
		);
//A5A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B9(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[324])
		);
//A5A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B10(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[325])
		);
//A5A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B11(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[326])
		);
//A5A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B12(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[327])
		);
//A5A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B13(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[328])
		);
//A5A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B14(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[329])
		);
//A5A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B15(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[330])
		);
//A5A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B16(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[331])
		);
//A5A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B17(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[332])
		);
//A5A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B18(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[333])
		);
//A5A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B19(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[334])
		);
//A5A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B20(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[335])
		);
//A5A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B21(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[336])
		);
//A5A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B22(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[337])
		);
//A5A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B23(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[338])
		);
//A5A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B24(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[339])
		);
//A5A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B25(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[340])
		);
//A5A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B26(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[341])
		);
//A5A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B27(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[342])
		);
//A5A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B28(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[343])
		);
//A5A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B29(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[344])
		);
//A5A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B30(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[345])
		);
//A5A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B31(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[346])
		);
//A5A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B32(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[347])
		);
//A5A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B33(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[348])
		);
//A5A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B34(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[349])
		);
//A5A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B35(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[350])
		);
//A5A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B36(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[351])
		);
//A5A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B37(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[352])
		);
//A5A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B38(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[353])
		);
//A5A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B39(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[354])
		);
//A5A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B40(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[355])
		);
//A5A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B41(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[356])
		);
//A5A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B42(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[357])
		);
//A5A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B43(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[358])
		);
//A5A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B44(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[359])
		);
//A5A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B45(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[360])
		);
//A5A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B46(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[361])
		);
//A5A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B47(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[362])
		);
//A5A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B48(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[363])
		);
//A5A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B49(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[364])
		);
//A5A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B50(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[365])
		);
//A5A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B51(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[366])
		);
//A5A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B52(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[367])
		);
//A5A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B53(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[368])
		);
//A5A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B54(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[369])
		);
//A5A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B55(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[370])
		);
//A5A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B56(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[371])
		);
//A5A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B57(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[372])
		);
//A5A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B58(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[373])
		);
//A5A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B59(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[374])
		);
//A5A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B60(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[375])
		);
//A5A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B61(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[376])
		);
//A5A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B62(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[377])
		);
//A5A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B63(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[378])
		);
//A5A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B64(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[379])
		);
//A5A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A5B65(
		.clk(clk),
			.A(A[5][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[380])
		);
//A6A6
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B6(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[6][BIT_LEN-1:0]),
			.P(mul_result[381])
		);
//A6A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B7(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[382])
		);
//A6A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B8(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[383])
		);
//A6A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B9(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[384])
		);
//A6A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B10(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[385])
		);
//A6A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B11(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[386])
		);
//A6A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B12(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[387])
		);
//A6A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B13(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[388])
		);
//A6A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B14(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[389])
		);
//A6A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B15(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[390])
		);
//A6A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B16(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[391])
		);
//A6A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B17(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[392])
		);
//A6A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B18(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[393])
		);
//A6A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B19(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[394])
		);
//A6A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B20(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[395])
		);
//A6A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B21(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[396])
		);
//A6A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B22(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[397])
		);
//A6A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B23(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[398])
		);
//A6A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B24(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[399])
		);
//A6A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B25(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[400])
		);
//A6A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B26(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[401])
		);
//A6A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B27(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[402])
		);
//A6A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B28(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[403])
		);
//A6A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B29(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[404])
		);
//A6A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B30(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[405])
		);
//A6A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B31(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[406])
		);
//A6A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B32(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[407])
		);
//A6A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B33(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[408])
		);
//A6A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B34(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[409])
		);
//A6A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B35(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[410])
		);
//A6A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B36(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[411])
		);
//A6A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B37(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[412])
		);
//A6A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B38(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[413])
		);
//A6A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B39(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[414])
		);
//A6A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B40(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[415])
		);
//A6A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B41(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[416])
		);
//A6A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B42(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[417])
		);
//A6A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B43(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[418])
		);
//A6A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B44(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[419])
		);
//A6A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B45(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[420])
		);
//A6A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B46(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[421])
		);
//A6A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B47(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[422])
		);
//A6A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B48(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[423])
		);
//A6A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B49(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[424])
		);
//A6A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B50(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[425])
		);
//A6A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B51(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[426])
		);
//A6A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B52(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[427])
		);
//A6A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B53(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[428])
		);
//A6A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B54(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[429])
		);
//A6A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B55(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[430])
		);
//A6A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B56(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[431])
		);
//A6A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B57(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[432])
		);
//A6A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B58(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[433])
		);
//A6A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B59(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[434])
		);
//A6A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B60(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[435])
		);
//A6A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B61(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[436])
		);
//A6A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B62(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[437])
		);
//A6A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B63(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[438])
		);
//A6A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B64(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[439])
		);
//A6A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A6B65(
		.clk(clk),
			.A(A[6][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[440])
		);
//A7A7
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B7(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[7][BIT_LEN-1:0]),
			.P(mul_result[441])
		);
//A7A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B8(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[442])
		);
//A7A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B9(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[443])
		);
//A7A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B10(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[444])
		);
//A7A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B11(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[445])
		);
//A7A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B12(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[446])
		);
//A7A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B13(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[447])
		);
//A7A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B14(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[448])
		);
//A7A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B15(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[449])
		);
//A7A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B16(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[450])
		);
//A7A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B17(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[451])
		);
//A7A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B18(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[452])
		);
//A7A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B19(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[453])
		);
//A7A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B20(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[454])
		);
//A7A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B21(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[455])
		);
//A7A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B22(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[456])
		);
//A7A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B23(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[457])
		);
//A7A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B24(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[458])
		);
//A7A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B25(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[459])
		);
//A7A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B26(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[460])
		);
//A7A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B27(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[461])
		);
//A7A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B28(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[462])
		);
//A7A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B29(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[463])
		);
//A7A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B30(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[464])
		);
//A7A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B31(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[465])
		);
//A7A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B32(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[466])
		);
//A7A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B33(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[467])
		);
//A7A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B34(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[468])
		);
//A7A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B35(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[469])
		);
//A7A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B36(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[470])
		);
//A7A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B37(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[471])
		);
//A7A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B38(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[472])
		);
//A7A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B39(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[473])
		);
//A7A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B40(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[474])
		);
//A7A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B41(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[475])
		);
//A7A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B42(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[476])
		);
//A7A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B43(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[477])
		);
//A7A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B44(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[478])
		);
//A7A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B45(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[479])
		);
//A7A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B46(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[480])
		);
//A7A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B47(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[481])
		);
//A7A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B48(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[482])
		);
//A7A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B49(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[483])
		);
//A7A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B50(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[484])
		);
//A7A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B51(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[485])
		);
//A7A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B52(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[486])
		);
//A7A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B53(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[487])
		);
//A7A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B54(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[488])
		);
//A7A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B55(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[489])
		);
//A7A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B56(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[490])
		);
//A7A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B57(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[491])
		);
//A7A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B58(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[492])
		);
//A7A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B59(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[493])
		);
//A7A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B60(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[494])
		);
//A7A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B61(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[495])
		);
//A7A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B62(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[496])
		);
//A7A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B63(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[497])
		);
//A7A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B64(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[498])
		);
//A7A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A7B65(
		.clk(clk),
			.A(A[7][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[499])
		);
//A8A8
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B8(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[8][BIT_LEN-1:0]),
			.P(mul_result[500])
		);
//A8A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B9(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[501])
		);
//A8A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B10(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[502])
		);
//A8A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B11(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[503])
		);
//A8A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B12(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[504])
		);
//A8A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B13(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[505])
		);
//A8A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B14(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[506])
		);
//A8A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B15(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[507])
		);
//A8A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B16(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[508])
		);
//A8A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B17(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[509])
		);
//A8A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B18(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[510])
		);
//A8A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B19(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[511])
		);
//A8A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B20(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[512])
		);
//A8A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B21(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[513])
		);
//A8A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B22(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[514])
		);
//A8A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B23(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[515])
		);
//A8A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B24(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[516])
		);
//A8A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B25(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[517])
		);
//A8A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B26(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[518])
		);
//A8A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B27(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[519])
		);
//A8A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B28(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[520])
		);
//A8A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B29(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[521])
		);
//A8A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B30(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[522])
		);
//A8A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B31(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[523])
		);
//A8A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B32(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[524])
		);
//A8A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B33(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[525])
		);
//A8A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B34(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[526])
		);
//A8A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B35(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[527])
		);
//A8A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B36(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[528])
		);
//A8A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B37(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[529])
		);
//A8A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B38(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[530])
		);
//A8A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B39(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[531])
		);
//A8A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B40(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[532])
		);
//A8A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B41(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[533])
		);
//A8A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B42(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[534])
		);
//A8A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B43(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[535])
		);
//A8A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B44(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[536])
		);
//A8A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B45(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[537])
		);
//A8A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B46(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[538])
		);
//A8A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B47(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[539])
		);
//A8A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B48(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[540])
		);
//A8A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B49(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[541])
		);
//A8A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B50(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[542])
		);
//A8A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B51(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[543])
		);
//A8A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B52(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[544])
		);
//A8A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B53(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[545])
		);
//A8A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B54(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[546])
		);
//A8A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B55(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[547])
		);
//A8A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B56(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[548])
		);
//A8A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B57(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[549])
		);
//A8A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B58(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[550])
		);
//A8A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B59(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[551])
		);
//A8A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B60(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[552])
		);
//A8A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B61(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[553])
		);
//A8A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B62(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[554])
		);
//A8A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B63(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[555])
		);
//A8A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B64(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[556])
		);
//A8A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A8B65(
		.clk(clk),
			.A(A[8][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[557])
		);
//A9A9
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B9(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[9][BIT_LEN-1:0]),
			.P(mul_result[558])
		);
//A9A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B10(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[559])
		);
//A9A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B11(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[560])
		);
//A9A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B12(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[561])
		);
//A9A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B13(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[562])
		);
//A9A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B14(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[563])
		);
//A9A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B15(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[564])
		);
//A9A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B16(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[565])
		);
//A9A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B17(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[566])
		);
//A9A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B18(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[567])
		);
//A9A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B19(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[568])
		);
//A9A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B20(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[569])
		);
//A9A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B21(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[570])
		);
//A9A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B22(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[571])
		);
//A9A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B23(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[572])
		);
//A9A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B24(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[573])
		);
//A9A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B25(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[574])
		);
//A9A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B26(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[575])
		);
//A9A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B27(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[576])
		);
//A9A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B28(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[577])
		);
//A9A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B29(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[578])
		);
//A9A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B30(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[579])
		);
//A9A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B31(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[580])
		);
//A9A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B32(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[581])
		);
//A9A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B33(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[582])
		);
//A9A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B34(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[583])
		);
//A9A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B35(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[584])
		);
//A9A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B36(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[585])
		);
//A9A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B37(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[586])
		);
//A9A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B38(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[587])
		);
//A9A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B39(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[588])
		);
//A9A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B40(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[589])
		);
//A9A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B41(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[590])
		);
//A9A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B42(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[591])
		);
//A9A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B43(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[592])
		);
//A9A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B44(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[593])
		);
//A9A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B45(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[594])
		);
//A9A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B46(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[595])
		);
//A9A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B47(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[596])
		);
//A9A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B48(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[597])
		);
//A9A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B49(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[598])
		);
//A9A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B50(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[599])
		);
//A9A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B51(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[600])
		);
//A9A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B52(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[601])
		);
//A9A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B53(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[602])
		);
//A9A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B54(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[603])
		);
//A9A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B55(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[604])
		);
//A9A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B56(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[605])
		);
//A9A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B57(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[606])
		);
//A9A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B58(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[607])
		);
//A9A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B59(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[608])
		);
//A9A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B60(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[609])
		);
//A9A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B61(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[610])
		);
//A9A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B62(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[611])
		);
//A9A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B63(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[612])
		);
//A9A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B64(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[613])
		);
//A9A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A9B65(
		.clk(clk),
			.A(A[9][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[614])
		);
//A10A10
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B10(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[10][BIT_LEN-1:0]),
			.P(mul_result[615])
		);
//A10A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B11(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[616])
		);
//A10A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B12(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[617])
		);
//A10A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B13(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[618])
		);
//A10A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B14(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[619])
		);
//A10A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B15(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[620])
		);
//A10A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B16(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[621])
		);
//A10A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B17(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[622])
		);
//A10A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B18(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[623])
		);
//A10A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B19(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[624])
		);
//A10A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B20(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[625])
		);
//A10A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B21(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[626])
		);
//A10A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B22(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[627])
		);
//A10A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B23(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[628])
		);
//A10A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B24(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[629])
		);
//A10A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B25(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[630])
		);
//A10A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B26(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[631])
		);
//A10A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B27(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[632])
		);
//A10A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B28(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[633])
		);
//A10A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B29(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[634])
		);
//A10A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B30(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[635])
		);
//A10A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B31(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[636])
		);
//A10A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B32(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[637])
		);
//A10A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B33(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[638])
		);
//A10A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B34(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[639])
		);
//A10A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B35(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[640])
		);
//A10A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B36(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[641])
		);
//A10A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B37(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[642])
		);
//A10A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B38(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[643])
		);
//A10A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B39(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[644])
		);
//A10A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B40(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[645])
		);
//A10A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B41(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[646])
		);
//A10A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B42(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[647])
		);
//A10A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B43(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[648])
		);
//A10A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B44(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[649])
		);
//A10A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B45(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[650])
		);
//A10A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B46(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[651])
		);
//A10A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B47(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[652])
		);
//A10A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B48(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[653])
		);
//A10A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B49(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[654])
		);
//A10A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B50(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[655])
		);
//A10A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B51(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[656])
		);
//A10A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B52(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[657])
		);
//A10A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B53(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[658])
		);
//A10A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B54(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[659])
		);
//A10A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B55(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[660])
		);
//A10A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B56(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[661])
		);
//A10A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B57(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[662])
		);
//A10A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B58(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[663])
		);
//A10A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B59(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[664])
		);
//A10A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B60(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[665])
		);
//A10A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B61(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[666])
		);
//A10A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B62(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[667])
		);
//A10A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B63(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[668])
		);
//A10A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B64(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[669])
		);
//A10A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A10B65(
		.clk(clk),
			.A(A[10][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[670])
		);
//A11A11
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B11(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[11][BIT_LEN-1:0]),
			.P(mul_result[671])
		);
//A11A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B12(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[672])
		);
//A11A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B13(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[673])
		);
//A11A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B14(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[674])
		);
//A11A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B15(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[675])
		);
//A11A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B16(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[676])
		);
//A11A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B17(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[677])
		);
//A11A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B18(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[678])
		);
//A11A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B19(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[679])
		);
//A11A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B20(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[680])
		);
//A11A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B21(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[681])
		);
//A11A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B22(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[682])
		);
//A11A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B23(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[683])
		);
//A11A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B24(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[684])
		);
//A11A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B25(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[685])
		);
//A11A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B26(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[686])
		);
//A11A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B27(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[687])
		);
//A11A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B28(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[688])
		);
//A11A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B29(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[689])
		);
//A11A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B30(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[690])
		);
//A11A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B31(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[691])
		);
//A11A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B32(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[692])
		);
//A11A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B33(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[693])
		);
//A11A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B34(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[694])
		);
//A11A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B35(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[695])
		);
//A11A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B36(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[696])
		);
//A11A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B37(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[697])
		);
//A11A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B38(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[698])
		);
//A11A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B39(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[699])
		);
//A11A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B40(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[700])
		);
//A11A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B41(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[701])
		);
//A11A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B42(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[702])
		);
//A11A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B43(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[703])
		);
//A11A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B44(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[704])
		);
//A11A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B45(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[705])
		);
//A11A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B46(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[706])
		);
//A11A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B47(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[707])
		);
//A11A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B48(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[708])
		);
//A11A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B49(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[709])
		);
//A11A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B50(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[710])
		);
//A11A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B51(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[711])
		);
//A11A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B52(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[712])
		);
//A11A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B53(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[713])
		);
//A11A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B54(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[714])
		);
//A11A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B55(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[715])
		);
//A11A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B56(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[716])
		);
//A11A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B57(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[717])
		);
//A11A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B58(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[718])
		);
//A11A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B59(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[719])
		);
//A11A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B60(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[720])
		);
//A11A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B61(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[721])
		);
//A11A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B62(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[722])
		);
//A11A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B63(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[723])
		);
//A11A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B64(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[724])
		);
//A11A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A11B65(
		.clk(clk),
			.A(A[11][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[725])
		);
//A12A12
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B12(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[12][BIT_LEN-1:0]),
			.P(mul_result[726])
		);
//A12A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B13(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[727])
		);
//A12A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B14(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[728])
		);
//A12A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B15(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[729])
		);
//A12A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B16(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[730])
		);
//A12A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B17(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[731])
		);
//A12A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B18(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[732])
		);
//A12A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B19(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[733])
		);
//A12A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B20(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[734])
		);
//A12A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B21(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[735])
		);
//A12A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B22(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[736])
		);
//A12A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B23(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[737])
		);
//A12A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B24(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[738])
		);
//A12A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B25(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[739])
		);
//A12A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B26(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[740])
		);
//A12A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B27(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[741])
		);
//A12A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B28(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[742])
		);
//A12A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B29(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[743])
		);
//A12A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B30(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[744])
		);
//A12A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B31(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[745])
		);
//A12A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B32(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[746])
		);
//A12A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B33(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[747])
		);
//A12A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B34(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[748])
		);
//A12A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B35(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[749])
		);
//A12A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B36(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[750])
		);
//A12A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B37(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[751])
		);
//A12A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B38(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[752])
		);
//A12A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B39(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[753])
		);
//A12A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B40(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[754])
		);
//A12A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B41(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[755])
		);
//A12A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B42(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[756])
		);
//A12A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B43(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[757])
		);
//A12A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B44(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[758])
		);
//A12A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B45(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[759])
		);
//A12A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B46(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[760])
		);
//A12A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B47(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[761])
		);
//A12A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B48(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[762])
		);
//A12A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B49(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[763])
		);
//A12A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B50(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[764])
		);
//A12A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B51(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[765])
		);
//A12A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B52(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[766])
		);
//A12A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B53(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[767])
		);
//A12A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B54(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[768])
		);
//A12A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B55(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[769])
		);
//A12A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B56(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[770])
		);
//A12A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B57(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[771])
		);
//A12A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B58(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[772])
		);
//A12A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B59(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[773])
		);
//A12A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B60(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[774])
		);
//A12A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B61(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[775])
		);
//A12A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B62(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[776])
		);
//A12A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B63(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[777])
		);
//A12A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B64(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[778])
		);
//A12A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A12B65(
		.clk(clk),
			.A(A[12][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[779])
		);
//A13A13
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B13(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[13][BIT_LEN-1:0]),
			.P(mul_result[780])
		);
//A13A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B14(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[781])
		);
//A13A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B15(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[782])
		);
//A13A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B16(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[783])
		);
//A13A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B17(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[784])
		);
//A13A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B18(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[785])
		);
//A13A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B19(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[786])
		);
//A13A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B20(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[787])
		);
//A13A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B21(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[788])
		);
//A13A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B22(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[789])
		);
//A13A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B23(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[790])
		);
//A13A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B24(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[791])
		);
//A13A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B25(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[792])
		);
//A13A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B26(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[793])
		);
//A13A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B27(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[794])
		);
//A13A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B28(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[795])
		);
//A13A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B29(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[796])
		);
//A13A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B30(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[797])
		);
//A13A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B31(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[798])
		);
//A13A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B32(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[799])
		);
//A13A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B33(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[800])
		);
//A13A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B34(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[801])
		);
//A13A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B35(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[802])
		);
//A13A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B36(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[803])
		);
//A13A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B37(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[804])
		);
//A13A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B38(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[805])
		);
//A13A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B39(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[806])
		);
//A13A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B40(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[807])
		);
//A13A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B41(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[808])
		);
//A13A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B42(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[809])
		);
//A13A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B43(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[810])
		);
//A13A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B44(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[811])
		);
//A13A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B45(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[812])
		);
//A13A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B46(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[813])
		);
//A13A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B47(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[814])
		);
//A13A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B48(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[815])
		);
//A13A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B49(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[816])
		);
//A13A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B50(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[817])
		);
//A13A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B51(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[818])
		);
//A13A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B52(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[819])
		);
//A13A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B53(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[820])
		);
//A13A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B54(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[821])
		);
//A13A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B55(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[822])
		);
//A13A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B56(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[823])
		);
//A13A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B57(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[824])
		);
//A13A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B58(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[825])
		);
//A13A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B59(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[826])
		);
//A13A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B60(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[827])
		);
//A13A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B61(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[828])
		);
//A13A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B62(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[829])
		);
//A13A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B63(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[830])
		);
//A13A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B64(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[831])
		);
//A13A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A13B65(
		.clk(clk),
			.A(A[13][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[832])
		);
//A14A14
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B14(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[14][BIT_LEN-1:0]),
			.P(mul_result[833])
		);
//A14A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B15(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[834])
		);
//A14A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B16(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[835])
		);
//A14A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B17(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[836])
		);
//A14A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B18(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[837])
		);
//A14A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B19(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[838])
		);
//A14A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B20(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[839])
		);
//A14A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B21(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[840])
		);
//A14A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B22(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[841])
		);
//A14A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B23(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[842])
		);
//A14A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B24(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[843])
		);
//A14A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B25(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[844])
		);
//A14A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B26(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[845])
		);
//A14A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B27(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[846])
		);
//A14A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B28(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[847])
		);
//A14A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B29(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[848])
		);
//A14A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B30(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[849])
		);
//A14A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B31(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[850])
		);
//A14A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B32(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[851])
		);
//A14A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B33(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[852])
		);
//A14A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B34(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[853])
		);
//A14A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B35(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[854])
		);
//A14A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B36(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[855])
		);
//A14A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B37(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[856])
		);
//A14A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B38(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[857])
		);
//A14A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B39(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[858])
		);
//A14A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B40(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[859])
		);
//A14A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B41(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[860])
		);
//A14A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B42(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[861])
		);
//A14A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B43(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[862])
		);
//A14A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B44(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[863])
		);
//A14A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B45(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[864])
		);
//A14A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B46(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[865])
		);
//A14A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B47(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[866])
		);
//A14A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B48(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[867])
		);
//A14A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B49(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[868])
		);
//A14A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B50(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[869])
		);
//A14A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B51(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[870])
		);
//A14A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B52(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[871])
		);
//A14A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B53(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[872])
		);
//A14A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B54(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[873])
		);
//A14A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B55(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[874])
		);
//A14A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B56(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[875])
		);
//A14A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B57(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[876])
		);
//A14A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B58(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[877])
		);
//A14A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B59(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[878])
		);
//A14A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B60(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[879])
		);
//A14A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B61(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[880])
		);
//A14A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B62(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[881])
		);
//A14A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B63(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[882])
		);
//A14A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B64(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[883])
		);
//A14A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A14B65(
		.clk(clk),
			.A(A[14][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[884])
		);
//A15A15
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B15(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[15][BIT_LEN-1:0]),
			.P(mul_result[885])
		);
//A15A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B16(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[886])
		);
//A15A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B17(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[887])
		);
//A15A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B18(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[888])
		);
//A15A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B19(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[889])
		);
//A15A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B20(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[890])
		);
//A15A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B21(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[891])
		);
//A15A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B22(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[892])
		);
//A15A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B23(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[893])
		);
//A15A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B24(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[894])
		);
//A15A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B25(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[895])
		);
//A15A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B26(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[896])
		);
//A15A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B27(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[897])
		);
//A15A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B28(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[898])
		);
//A15A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B29(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[899])
		);
//A15A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B30(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[900])
		);
//A15A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B31(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[901])
		);
//A15A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B32(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[902])
		);
//A15A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B33(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[903])
		);
//A15A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B34(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[904])
		);
//A15A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B35(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[905])
		);
//A15A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B36(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[906])
		);
//A15A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B37(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[907])
		);
//A15A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B38(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[908])
		);
//A15A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B39(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[909])
		);
//A15A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B40(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[910])
		);
//A15A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B41(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[911])
		);
//A15A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B42(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[912])
		);
//A15A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B43(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[913])
		);
//A15A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B44(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[914])
		);
//A15A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B45(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[915])
		);
//A15A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B46(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[916])
		);
//A15A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B47(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[917])
		);
//A15A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B48(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[918])
		);
//A15A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B49(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[919])
		);
//A15A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B50(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[920])
		);
//A15A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B51(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[921])
		);
//A15A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B52(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[922])
		);
//A15A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B53(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[923])
		);
//A15A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B54(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[924])
		);
//A15A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B55(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[925])
		);
//A15A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B56(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[926])
		);
//A15A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B57(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[927])
		);
//A15A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B58(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[928])
		);
//A15A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B59(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[929])
		);
//A15A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B60(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[930])
		);
//A15A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B61(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[931])
		);
//A15A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B62(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[932])
		);
//A15A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B63(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[933])
		);
//A15A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B64(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[934])
		);
//A15A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A15B65(
		.clk(clk),
			.A(A[15][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[935])
		);
//A16A16
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B16(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[16][BIT_LEN-1:0]),
			.P(mul_result[936])
		);
//A16A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B17(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[937])
		);
//A16A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B18(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[938])
		);
//A16A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B19(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[939])
		);
//A16A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B20(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[940])
		);
//A16A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B21(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[941])
		);
//A16A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B22(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[942])
		);
//A16A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B23(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[943])
		);
//A16A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B24(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[944])
		);
//A16A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B25(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[945])
		);
//A16A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B26(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[946])
		);
//A16A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B27(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[947])
		);
//A16A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B28(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[948])
		);
//A16A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B29(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[949])
		);
//A16A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B30(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[950])
		);
//A16A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B31(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[951])
		);
//A16A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B32(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[952])
		);
//A16A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B33(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[953])
		);
//A16A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B34(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[954])
		);
//A16A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B35(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[955])
		);
//A16A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B36(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[956])
		);
//A16A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B37(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[957])
		);
//A16A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B38(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[958])
		);
//A16A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B39(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[959])
		);
//A16A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B40(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[960])
		);
//A16A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B41(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[961])
		);
//A16A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B42(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[962])
		);
//A16A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B43(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[963])
		);
//A16A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B44(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[964])
		);
//A16A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B45(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[965])
		);
//A16A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B46(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[966])
		);
//A16A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B47(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[967])
		);
//A16A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B48(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[968])
		);
//A16A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B49(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[969])
		);
//A16A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B50(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[970])
		);
//A16A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B51(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[971])
		);
//A16A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B52(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[972])
		);
//A16A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B53(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[973])
		);
//A16A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B54(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[974])
		);
//A16A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B55(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[975])
		);
//A16A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B56(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[976])
		);
//A16A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B57(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[977])
		);
//A16A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B58(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[978])
		);
//A16A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B59(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[979])
		);
//A16A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B60(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[980])
		);
//A16A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B61(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[981])
		);
//A16A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B62(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[982])
		);
//A16A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B63(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[983])
		);
//A16A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B64(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[984])
		);
//A16A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A16B65(
		.clk(clk),
			.A(A[16][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[985])
		);
//A17A17
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B17(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[17][BIT_LEN-1:0]),
			.P(mul_result[986])
		);
//A17A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B18(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[987])
		);
//A17A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B19(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[988])
		);
//A17A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B20(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[989])
		);
//A17A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B21(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[990])
		);
//A17A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B22(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[991])
		);
//A17A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B23(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[992])
		);
//A17A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B24(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[993])
		);
//A17A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B25(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[994])
		);
//A17A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B26(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[995])
		);
//A17A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B27(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[996])
		);
//A17A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B28(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[997])
		);
//A17A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B29(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[998])
		);
//A17A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B30(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[999])
		);
//A17A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B31(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1000])
		);
//A17A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B32(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1001])
		);
//A17A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B33(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1002])
		);
//A17A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B34(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1003])
		);
//A17A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B35(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1004])
		);
//A17A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B36(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1005])
		);
//A17A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B37(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1006])
		);
//A17A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B38(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1007])
		);
//A17A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B39(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1008])
		);
//A17A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B40(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1009])
		);
//A17A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B41(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1010])
		);
//A17A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B42(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1011])
		);
//A17A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B43(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1012])
		);
//A17A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B44(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1013])
		);
//A17A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B45(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1014])
		);
//A17A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B46(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1015])
		);
//A17A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B47(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1016])
		);
//A17A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B48(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1017])
		);
//A17A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B49(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1018])
		);
//A17A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B50(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1019])
		);
//A17A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B51(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1020])
		);
//A17A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B52(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1021])
		);
//A17A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B53(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1022])
		);
//A17A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B54(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1023])
		);
//A17A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B55(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1024])
		);
//A17A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B56(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1025])
		);
//A17A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B57(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1026])
		);
//A17A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B58(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1027])
		);
//A17A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B59(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1028])
		);
//A17A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B60(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1029])
		);
//A17A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B61(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1030])
		);
//A17A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B62(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1031])
		);
//A17A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B63(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1032])
		);
//A17A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B64(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1033])
		);
//A17A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A17B65(
		.clk(clk),
			.A(A[17][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1034])
		);
//A18A18
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B18(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[18][BIT_LEN-1:0]),
			.P(mul_result[1035])
		);
//A18A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B19(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[1036])
		);
//A18A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B20(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[1037])
		);
//A18A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B21(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[1038])
		);
//A18A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B22(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[1039])
		);
//A18A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B23(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[1040])
		);
//A18A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B24(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[1041])
		);
//A18A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B25(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1042])
		);
//A18A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B26(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1043])
		);
//A18A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B27(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1044])
		);
//A18A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B28(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1045])
		);
//A18A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B29(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1046])
		);
//A18A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B30(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1047])
		);
//A18A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B31(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1048])
		);
//A18A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B32(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1049])
		);
//A18A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B33(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1050])
		);
//A18A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B34(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1051])
		);
//A18A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B35(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1052])
		);
//A18A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B36(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1053])
		);
//A18A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B37(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1054])
		);
//A18A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B38(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1055])
		);
//A18A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B39(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1056])
		);
//A18A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B40(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1057])
		);
//A18A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B41(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1058])
		);
//A18A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B42(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1059])
		);
//A18A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B43(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1060])
		);
//A18A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B44(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1061])
		);
//A18A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B45(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1062])
		);
//A18A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B46(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1063])
		);
//A18A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B47(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1064])
		);
//A18A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B48(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1065])
		);
//A18A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B49(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1066])
		);
//A18A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B50(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1067])
		);
//A18A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B51(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1068])
		);
//A18A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B52(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1069])
		);
//A18A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B53(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1070])
		);
//A18A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B54(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1071])
		);
//A18A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B55(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1072])
		);
//A18A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B56(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1073])
		);
//A18A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B57(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1074])
		);
//A18A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B58(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1075])
		);
//A18A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B59(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1076])
		);
//A18A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B60(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1077])
		);
//A18A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B61(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1078])
		);
//A18A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B62(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1079])
		);
//A18A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B63(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1080])
		);
//A18A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B64(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1081])
		);
//A18A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A18B65(
		.clk(clk),
			.A(A[18][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1082])
		);
//A19A19
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B19(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[19][BIT_LEN-1:0]),
			.P(mul_result[1083])
		);
//A19A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B20(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[1084])
		);
//A19A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B21(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[1085])
		);
//A19A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B22(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[1086])
		);
//A19A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B23(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[1087])
		);
//A19A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B24(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[1088])
		);
//A19A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B25(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1089])
		);
//A19A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B26(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1090])
		);
//A19A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B27(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1091])
		);
//A19A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B28(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1092])
		);
//A19A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B29(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1093])
		);
//A19A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B30(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1094])
		);
//A19A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B31(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1095])
		);
//A19A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B32(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1096])
		);
//A19A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B33(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1097])
		);
//A19A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B34(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1098])
		);
//A19A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B35(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1099])
		);
//A19A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B36(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1100])
		);
//A19A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B37(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1101])
		);
//A19A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B38(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1102])
		);
//A19A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B39(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1103])
		);
//A19A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B40(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1104])
		);
//A19A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B41(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1105])
		);
//A19A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B42(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1106])
		);
//A19A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B43(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1107])
		);
//A19A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B44(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1108])
		);
//A19A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B45(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1109])
		);
//A19A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B46(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1110])
		);
//A19A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B47(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1111])
		);
//A19A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B48(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1112])
		);
//A19A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B49(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1113])
		);
//A19A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B50(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1114])
		);
//A19A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B51(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1115])
		);
//A19A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B52(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1116])
		);
//A19A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B53(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1117])
		);
//A19A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B54(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1118])
		);
//A19A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B55(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1119])
		);
//A19A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B56(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1120])
		);
//A19A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B57(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1121])
		);
//A19A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B58(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1122])
		);
//A19A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B59(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1123])
		);
//A19A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B60(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1124])
		);
//A19A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B61(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1125])
		);
//A19A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B62(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1126])
		);
//A19A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B63(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1127])
		);
//A19A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B64(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1128])
		);
//A19A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A19B65(
		.clk(clk),
			.A(A[19][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1129])
		);
//A20A20
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B20(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[20][BIT_LEN-1:0]),
			.P(mul_result[1130])
		);
//A20A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B21(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[1131])
		);
//A20A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B22(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[1132])
		);
//A20A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B23(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[1133])
		);
//A20A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B24(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[1134])
		);
//A20A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B25(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1135])
		);
//A20A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B26(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1136])
		);
//A20A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B27(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1137])
		);
//A20A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B28(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1138])
		);
//A20A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B29(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1139])
		);
//A20A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B30(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1140])
		);
//A20A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B31(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1141])
		);
//A20A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B32(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1142])
		);
//A20A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B33(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1143])
		);
//A20A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B34(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1144])
		);
//A20A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B35(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1145])
		);
//A20A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B36(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1146])
		);
//A20A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B37(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1147])
		);
//A20A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B38(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1148])
		);
//A20A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B39(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1149])
		);
//A20A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B40(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1150])
		);
//A20A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B41(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1151])
		);
//A20A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B42(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1152])
		);
//A20A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B43(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1153])
		);
//A20A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B44(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1154])
		);
//A20A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B45(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1155])
		);
//A20A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B46(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1156])
		);
//A20A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B47(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1157])
		);
//A20A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B48(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1158])
		);
//A20A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B49(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1159])
		);
//A20A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B50(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1160])
		);
//A20A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B51(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1161])
		);
//A20A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B52(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1162])
		);
//A20A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B53(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1163])
		);
//A20A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B54(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1164])
		);
//A20A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B55(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1165])
		);
//A20A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B56(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1166])
		);
//A20A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B57(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1167])
		);
//A20A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B58(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1168])
		);
//A20A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B59(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1169])
		);
//A20A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B60(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1170])
		);
//A20A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B61(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1171])
		);
//A20A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B62(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1172])
		);
//A20A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B63(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1173])
		);
//A20A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B64(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1174])
		);
//A20A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A20B65(
		.clk(clk),
			.A(A[20][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1175])
		);
//A21A21
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B21(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[21][BIT_LEN-1:0]),
			.P(mul_result[1176])
		);
//A21A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B22(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[1177])
		);
//A21A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B23(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[1178])
		);
//A21A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B24(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[1179])
		);
//A21A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B25(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1180])
		);
//A21A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B26(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1181])
		);
//A21A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B27(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1182])
		);
//A21A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B28(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1183])
		);
//A21A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B29(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1184])
		);
//A21A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B30(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1185])
		);
//A21A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B31(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1186])
		);
//A21A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B32(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1187])
		);
//A21A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B33(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1188])
		);
//A21A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B34(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1189])
		);
//A21A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B35(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1190])
		);
//A21A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B36(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1191])
		);
//A21A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B37(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1192])
		);
//A21A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B38(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1193])
		);
//A21A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B39(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1194])
		);
//A21A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B40(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1195])
		);
//A21A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B41(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1196])
		);
//A21A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B42(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1197])
		);
//A21A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B43(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1198])
		);
//A21A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B44(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1199])
		);
//A21A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B45(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1200])
		);
//A21A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B46(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1201])
		);
//A21A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B47(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1202])
		);
//A21A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B48(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1203])
		);
//A21A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B49(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1204])
		);
//A21A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B50(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1205])
		);
//A21A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B51(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1206])
		);
//A21A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B52(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1207])
		);
//A21A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B53(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1208])
		);
//A21A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B54(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1209])
		);
//A21A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B55(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1210])
		);
//A21A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B56(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1211])
		);
//A21A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B57(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1212])
		);
//A21A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B58(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1213])
		);
//A21A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B59(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1214])
		);
//A21A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B60(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1215])
		);
//A21A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B61(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1216])
		);
//A21A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B62(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1217])
		);
//A21A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B63(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1218])
		);
//A21A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B64(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1219])
		);
//A21A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A21B65(
		.clk(clk),
			.A(A[21][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1220])
		);
//A22A22
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B22(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[22][BIT_LEN-1:0]),
			.P(mul_result[1221])
		);
//A22A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B23(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[1222])
		);
//A22A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B24(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[1223])
		);
//A22A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B25(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1224])
		);
//A22A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B26(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1225])
		);
//A22A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B27(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1226])
		);
//A22A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B28(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1227])
		);
//A22A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B29(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1228])
		);
//A22A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B30(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1229])
		);
//A22A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B31(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1230])
		);
//A22A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B32(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1231])
		);
//A22A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B33(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1232])
		);
//A22A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B34(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1233])
		);
//A22A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B35(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1234])
		);
//A22A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B36(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1235])
		);
//A22A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B37(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1236])
		);
//A22A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B38(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1237])
		);
//A22A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B39(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1238])
		);
//A22A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B40(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1239])
		);
//A22A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B41(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1240])
		);
//A22A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B42(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1241])
		);
//A22A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B43(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1242])
		);
//A22A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B44(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1243])
		);
//A22A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B45(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1244])
		);
//A22A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B46(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1245])
		);
//A22A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B47(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1246])
		);
//A22A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B48(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1247])
		);
//A22A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B49(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1248])
		);
//A22A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B50(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1249])
		);
//A22A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B51(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1250])
		);
//A22A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B52(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1251])
		);
//A22A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B53(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1252])
		);
//A22A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B54(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1253])
		);
//A22A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B55(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1254])
		);
//A22A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B56(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1255])
		);
//A22A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B57(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1256])
		);
//A22A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B58(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1257])
		);
//A22A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B59(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1258])
		);
//A22A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B60(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1259])
		);
//A22A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B61(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1260])
		);
//A22A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B62(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1261])
		);
//A22A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B63(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1262])
		);
//A22A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B64(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1263])
		);
//A22A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A22B65(
		.clk(clk),
			.A(A[22][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1264])
		);
//A23A23
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B23(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[23][BIT_LEN-1:0]),
			.P(mul_result[1265])
		);
//A23A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B24(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[1266])
		);
//A23A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B25(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1267])
		);
//A23A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B26(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1268])
		);
//A23A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B27(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1269])
		);
//A23A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B28(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1270])
		);
//A23A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B29(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1271])
		);
//A23A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B30(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1272])
		);
//A23A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B31(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1273])
		);
//A23A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B32(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1274])
		);
//A23A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B33(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1275])
		);
//A23A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B34(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1276])
		);
//A23A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B35(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1277])
		);
//A23A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B36(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1278])
		);
//A23A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B37(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1279])
		);
//A23A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B38(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1280])
		);
//A23A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B39(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1281])
		);
//A23A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B40(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1282])
		);
//A23A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B41(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1283])
		);
//A23A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B42(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1284])
		);
//A23A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B43(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1285])
		);
//A23A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B44(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1286])
		);
//A23A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B45(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1287])
		);
//A23A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B46(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1288])
		);
//A23A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B47(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1289])
		);
//A23A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B48(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1290])
		);
//A23A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B49(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1291])
		);
//A23A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B50(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1292])
		);
//A23A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B51(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1293])
		);
//A23A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B52(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1294])
		);
//A23A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B53(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1295])
		);
//A23A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B54(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1296])
		);
//A23A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B55(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1297])
		);
//A23A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B56(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1298])
		);
//A23A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B57(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1299])
		);
//A23A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B58(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1300])
		);
//A23A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B59(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1301])
		);
//A23A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B60(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1302])
		);
//A23A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B61(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1303])
		);
//A23A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B62(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1304])
		);
//A23A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B63(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1305])
		);
//A23A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B64(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1306])
		);
//A23A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A23B65(
		.clk(clk),
			.A(A[23][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1307])
		);
//A24A24
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B24(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[24][BIT_LEN-1:0]),
			.P(mul_result[1308])
		);
//A24A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B25(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1309])
		);
//A24A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B26(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1310])
		);
//A24A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B27(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1311])
		);
//A24A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B28(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1312])
		);
//A24A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B29(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1313])
		);
//A24A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B30(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1314])
		);
//A24A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B31(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1315])
		);
//A24A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B32(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1316])
		);
//A24A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B33(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1317])
		);
//A24A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B34(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1318])
		);
//A24A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B35(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1319])
		);
//A24A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B36(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1320])
		);
//A24A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B37(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1321])
		);
//A24A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B38(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1322])
		);
//A24A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B39(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1323])
		);
//A24A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B40(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1324])
		);
//A24A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B41(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1325])
		);
//A24A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B42(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1326])
		);
//A24A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B43(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1327])
		);
//A24A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B44(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1328])
		);
//A24A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B45(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1329])
		);
//A24A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B46(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1330])
		);
//A24A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B47(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1331])
		);
//A24A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B48(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1332])
		);
//A24A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B49(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1333])
		);
//A24A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B50(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1334])
		);
//A24A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B51(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1335])
		);
//A24A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B52(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1336])
		);
//A24A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B53(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1337])
		);
//A24A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B54(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1338])
		);
//A24A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B55(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1339])
		);
//A24A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B56(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1340])
		);
//A24A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B57(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1341])
		);
//A24A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B58(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1342])
		);
//A24A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B59(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1343])
		);
//A24A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B60(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1344])
		);
//A24A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B61(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1345])
		);
//A24A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B62(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1346])
		);
//A24A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B63(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1347])
		);
//A24A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B64(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1348])
		);
//A24A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A24B65(
		.clk(clk),
			.A(A[24][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1349])
		);
//A25A25
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B25(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[25][BIT_LEN-1:0]),
			.P(mul_result[1350])
		);
//A25A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B26(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1351])
		);
//A25A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B27(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1352])
		);
//A25A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B28(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1353])
		);
//A25A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B29(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1354])
		);
//A25A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B30(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1355])
		);
//A25A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B31(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1356])
		);
//A25A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B32(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1357])
		);
//A25A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B33(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1358])
		);
//A25A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B34(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1359])
		);
//A25A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B35(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1360])
		);
//A25A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B36(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1361])
		);
//A25A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B37(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1362])
		);
//A25A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B38(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1363])
		);
//A25A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B39(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1364])
		);
//A25A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B40(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1365])
		);
//A25A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B41(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1366])
		);
//A25A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B42(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1367])
		);
//A25A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B43(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1368])
		);
//A25A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B44(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1369])
		);
//A25A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B45(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1370])
		);
//A25A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B46(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1371])
		);
//A25A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B47(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1372])
		);
//A25A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B48(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1373])
		);
//A25A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B49(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1374])
		);
//A25A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B50(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1375])
		);
//A25A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B51(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1376])
		);
//A25A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B52(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1377])
		);
//A25A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B53(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1378])
		);
//A25A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B54(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1379])
		);
//A25A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B55(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1380])
		);
//A25A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B56(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1381])
		);
//A25A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B57(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1382])
		);
//A25A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B58(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1383])
		);
//A25A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B59(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1384])
		);
//A25A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B60(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1385])
		);
//A25A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B61(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1386])
		);
//A25A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B62(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1387])
		);
//A25A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B63(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1388])
		);
//A25A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B64(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1389])
		);
//A25A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A25B65(
		.clk(clk),
			.A(A[25][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1390])
		);
//A26A26
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B26(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[26][BIT_LEN-1:0]),
			.P(mul_result[1391])
		);
//A26A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B27(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1392])
		);
//A26A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B28(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1393])
		);
//A26A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B29(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1394])
		);
//A26A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B30(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1395])
		);
//A26A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B31(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1396])
		);
//A26A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B32(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1397])
		);
//A26A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B33(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1398])
		);
//A26A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B34(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1399])
		);
//A26A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B35(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1400])
		);
//A26A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B36(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1401])
		);
//A26A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B37(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1402])
		);
//A26A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B38(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1403])
		);
//A26A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B39(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1404])
		);
//A26A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B40(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1405])
		);
//A26A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B41(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1406])
		);
//A26A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B42(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1407])
		);
//A26A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B43(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1408])
		);
//A26A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B44(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1409])
		);
//A26A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B45(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1410])
		);
//A26A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B46(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1411])
		);
//A26A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B47(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1412])
		);
//A26A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B48(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1413])
		);
//A26A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B49(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1414])
		);
//A26A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B50(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1415])
		);
//A26A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B51(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1416])
		);
//A26A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B52(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1417])
		);
//A26A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B53(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1418])
		);
//A26A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B54(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1419])
		);
//A26A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B55(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1420])
		);
//A26A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B56(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1421])
		);
//A26A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B57(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1422])
		);
//A26A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B58(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1423])
		);
//A26A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B59(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1424])
		);
//A26A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B60(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1425])
		);
//A26A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B61(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1426])
		);
//A26A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B62(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1427])
		);
//A26A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B63(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1428])
		);
//A26A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B64(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1429])
		);
//A26A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A26B65(
		.clk(clk),
			.A(A[26][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1430])
		);
//A27A27
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B27(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[27][BIT_LEN-1:0]),
			.P(mul_result[1431])
		);
//A27A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B28(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1432])
		);
//A27A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B29(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1433])
		);
//A27A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B30(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1434])
		);
//A27A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B31(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1435])
		);
//A27A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B32(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1436])
		);
//A27A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B33(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1437])
		);
//A27A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B34(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1438])
		);
//A27A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B35(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1439])
		);
//A27A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B36(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1440])
		);
//A27A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B37(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1441])
		);
//A27A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B38(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1442])
		);
//A27A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B39(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1443])
		);
//A27A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B40(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1444])
		);
//A27A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B41(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1445])
		);
//A27A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B42(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1446])
		);
//A27A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B43(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1447])
		);
//A27A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B44(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1448])
		);
//A27A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B45(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1449])
		);
//A27A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B46(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1450])
		);
//A27A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B47(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1451])
		);
//A27A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B48(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1452])
		);
//A27A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B49(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1453])
		);
//A27A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B50(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1454])
		);
//A27A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B51(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1455])
		);
//A27A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B52(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1456])
		);
//A27A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B53(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1457])
		);
//A27A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B54(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1458])
		);
//A27A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B55(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1459])
		);
//A27A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B56(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1460])
		);
//A27A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B57(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1461])
		);
//A27A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B58(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1462])
		);
//A27A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B59(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1463])
		);
//A27A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B60(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1464])
		);
//A27A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B61(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1465])
		);
//A27A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B62(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1466])
		);
//A27A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B63(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1467])
		);
//A27A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B64(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1468])
		);
//A27A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A27B65(
		.clk(clk),
			.A(A[27][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1469])
		);
//A28A28
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B28(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[28][BIT_LEN-1:0]),
			.P(mul_result[1470])
		);
//A28A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B29(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1471])
		);
//A28A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B30(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1472])
		);
//A28A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B31(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1473])
		);
//A28A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B32(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1474])
		);
//A28A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B33(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1475])
		);
//A28A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B34(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1476])
		);
//A28A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B35(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1477])
		);
//A28A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B36(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1478])
		);
//A28A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B37(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1479])
		);
//A28A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B38(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1480])
		);
//A28A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B39(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1481])
		);
//A28A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B40(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1482])
		);
//A28A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B41(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1483])
		);
//A28A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B42(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1484])
		);
//A28A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B43(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1485])
		);
//A28A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B44(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1486])
		);
//A28A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B45(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1487])
		);
//A28A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B46(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1488])
		);
//A28A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B47(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1489])
		);
//A28A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B48(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1490])
		);
//A28A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B49(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1491])
		);
//A28A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B50(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1492])
		);
//A28A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B51(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1493])
		);
//A28A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B52(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1494])
		);
//A28A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B53(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1495])
		);
//A28A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B54(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1496])
		);
//A28A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B55(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1497])
		);
//A28A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B56(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1498])
		);
//A28A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B57(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1499])
		);
//A28A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B58(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1500])
		);
//A28A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B59(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1501])
		);
//A28A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B60(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1502])
		);
//A28A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B61(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1503])
		);
//A28A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B62(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1504])
		);
//A28A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B63(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1505])
		);
//A28A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B64(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1506])
		);
//A28A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A28B65(
		.clk(clk),
			.A(A[28][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1507])
		);
//A29A29
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B29(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[29][BIT_LEN-1:0]),
			.P(mul_result[1508])
		);
//A29A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B30(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1509])
		);
//A29A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B31(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1510])
		);
//A29A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B32(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1511])
		);
//A29A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B33(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1512])
		);
//A29A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B34(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1513])
		);
//A29A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B35(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1514])
		);
//A29A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B36(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1515])
		);
//A29A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B37(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1516])
		);
//A29A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B38(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1517])
		);
//A29A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B39(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1518])
		);
//A29A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B40(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1519])
		);
//A29A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B41(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1520])
		);
//A29A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B42(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1521])
		);
//A29A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B43(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1522])
		);
//A29A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B44(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1523])
		);
//A29A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B45(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1524])
		);
//A29A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B46(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1525])
		);
//A29A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B47(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1526])
		);
//A29A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B48(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1527])
		);
//A29A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B49(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1528])
		);
//A29A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B50(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1529])
		);
//A29A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B51(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1530])
		);
//A29A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B52(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1531])
		);
//A29A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B53(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1532])
		);
//A29A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B54(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1533])
		);
//A29A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B55(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1534])
		);
//A29A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B56(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1535])
		);
//A29A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B57(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1536])
		);
//A29A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B58(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1537])
		);
//A29A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B59(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1538])
		);
//A29A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B60(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1539])
		);
//A29A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B61(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1540])
		);
//A29A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B62(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1541])
		);
//A29A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B63(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1542])
		);
//A29A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B64(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1543])
		);
//A29A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A29B65(
		.clk(clk),
			.A(A[29][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1544])
		);
//A30A30
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B30(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[30][BIT_LEN-1:0]),
			.P(mul_result[1545])
		);
//A30A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B31(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1546])
		);
//A30A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B32(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1547])
		);
//A30A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B33(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1548])
		);
//A30A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B34(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1549])
		);
//A30A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B35(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1550])
		);
//A30A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B36(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1551])
		);
//A30A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B37(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1552])
		);
//A30A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B38(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1553])
		);
//A30A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B39(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1554])
		);
//A30A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B40(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1555])
		);
//A30A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B41(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1556])
		);
//A30A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B42(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1557])
		);
//A30A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B43(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1558])
		);
//A30A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B44(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1559])
		);
//A30A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B45(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1560])
		);
//A30A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B46(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1561])
		);
//A30A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B47(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1562])
		);
//A30A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B48(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1563])
		);
//A30A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B49(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1564])
		);
//A30A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B50(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1565])
		);
//A30A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B51(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1566])
		);
//A30A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B52(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1567])
		);
//A30A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B53(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1568])
		);
//A30A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B54(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1569])
		);
//A30A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B55(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1570])
		);
//A30A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B56(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1571])
		);
//A30A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B57(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1572])
		);
//A30A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B58(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1573])
		);
//A30A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B59(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1574])
		);
//A30A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B60(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1575])
		);
//A30A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B61(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1576])
		);
//A30A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B62(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1577])
		);
//A30A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B63(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1578])
		);
//A30A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B64(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1579])
		);
//A30A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A30B65(
		.clk(clk),
			.A(A[30][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1580])
		);
//A31A31
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B31(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[31][BIT_LEN-1:0]),
			.P(mul_result[1581])
		);
//A31A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B32(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1582])
		);
//A31A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B33(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1583])
		);
//A31A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B34(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1584])
		);
//A31A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B35(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1585])
		);
//A31A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B36(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1586])
		);
//A31A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B37(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1587])
		);
//A31A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B38(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1588])
		);
//A31A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B39(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1589])
		);
//A31A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B40(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1590])
		);
//A31A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B41(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1591])
		);
//A31A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B42(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1592])
		);
//A31A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B43(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1593])
		);
//A31A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B44(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1594])
		);
//A31A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B45(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1595])
		);
//A31A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B46(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1596])
		);
//A31A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B47(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1597])
		);
//A31A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B48(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1598])
		);
//A31A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B49(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1599])
		);
//A31A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B50(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1600])
		);
//A31A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B51(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1601])
		);
//A31A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B52(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1602])
		);
//A31A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B53(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1603])
		);
//A31A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B54(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1604])
		);
//A31A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B55(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1605])
		);
//A31A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B56(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1606])
		);
//A31A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B57(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1607])
		);
//A31A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B58(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1608])
		);
//A31A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B59(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1609])
		);
//A31A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B60(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1610])
		);
//A31A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B61(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1611])
		);
//A31A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B62(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1612])
		);
//A31A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B63(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1613])
		);
//A31A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B64(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1614])
		);
//A31A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A31B65(
		.clk(clk),
			.A(A[31][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1615])
		);
//A32A32
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B32(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[32][BIT_LEN-1:0]),
			.P(mul_result[1616])
		);
//A32A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B33(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1617])
		);
//A32A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B34(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1618])
		);
//A32A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B35(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1619])
		);
//A32A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B36(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1620])
		);
//A32A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B37(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1621])
		);
//A32A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B38(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1622])
		);
//A32A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B39(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1623])
		);
//A32A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B40(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1624])
		);
//A32A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B41(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1625])
		);
//A32A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B42(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1626])
		);
//A32A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B43(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1627])
		);
//A32A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B44(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1628])
		);
//A32A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B45(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1629])
		);
//A32A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B46(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1630])
		);
//A32A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B47(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1631])
		);
//A32A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B48(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1632])
		);
//A32A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B49(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1633])
		);
//A32A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B50(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1634])
		);
//A32A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B51(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1635])
		);
//A32A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B52(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1636])
		);
//A32A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B53(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1637])
		);
//A32A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B54(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1638])
		);
//A32A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B55(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1639])
		);
//A32A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B56(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1640])
		);
//A32A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B57(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1641])
		);
//A32A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B58(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1642])
		);
//A32A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B59(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1643])
		);
//A32A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B60(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1644])
		);
//A32A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B61(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1645])
		);
//A32A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B62(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1646])
		);
//A32A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B63(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1647])
		);
//A32A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B64(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1648])
		);
//A32A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A32B65(
		.clk(clk),
			.A(A[32][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1649])
		);
//A33A33
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B33(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[33][BIT_LEN-1:0]),
			.P(mul_result[1650])
		);
//A33A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B34(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1651])
		);
//A33A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B35(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1652])
		);
//A33A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B36(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1653])
		);
//A33A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B37(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1654])
		);
//A33A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B38(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1655])
		);
//A33A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B39(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1656])
		);
//A33A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B40(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1657])
		);
//A33A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B41(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1658])
		);
//A33A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B42(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1659])
		);
//A33A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B43(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1660])
		);
//A33A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B44(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1661])
		);
//A33A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B45(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1662])
		);
//A33A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B46(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1663])
		);
//A33A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B47(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1664])
		);
//A33A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B48(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1665])
		);
//A33A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B49(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1666])
		);
//A33A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B50(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1667])
		);
//A33A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B51(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1668])
		);
//A33A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B52(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1669])
		);
//A33A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B53(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1670])
		);
//A33A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B54(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1671])
		);
//A33A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B55(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1672])
		);
//A33A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B56(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1673])
		);
//A33A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B57(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1674])
		);
//A33A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B58(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1675])
		);
//A33A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B59(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1676])
		);
//A33A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B60(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1677])
		);
//A33A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B61(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1678])
		);
//A33A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B62(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1679])
		);
//A33A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B63(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1680])
		);
//A33A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B64(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1681])
		);
//A33A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A33B65(
		.clk(clk),
			.A(A[33][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1682])
		);
//A34A34
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B34(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[34][BIT_LEN-1:0]),
			.P(mul_result[1683])
		);
//A34A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B35(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1684])
		);
//A34A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B36(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1685])
		);
//A34A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B37(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1686])
		);
//A34A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B38(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1687])
		);
//A34A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B39(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1688])
		);
//A34A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B40(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1689])
		);
//A34A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B41(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1690])
		);
//A34A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B42(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1691])
		);
//A34A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B43(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1692])
		);
//A34A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B44(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1693])
		);
//A34A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B45(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1694])
		);
//A34A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B46(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1695])
		);
//A34A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B47(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1696])
		);
//A34A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B48(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1697])
		);
//A34A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B49(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1698])
		);
//A34A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B50(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1699])
		);
//A34A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B51(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1700])
		);
//A34A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B52(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1701])
		);
//A34A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B53(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1702])
		);
//A34A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B54(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1703])
		);
//A34A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B55(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1704])
		);
//A34A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B56(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1705])
		);
//A34A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B57(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1706])
		);
//A34A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B58(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1707])
		);
//A34A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B59(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1708])
		);
//A34A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B60(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1709])
		);
//A34A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B61(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1710])
		);
//A34A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B62(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1711])
		);
//A34A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B63(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1712])
		);
//A34A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B64(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1713])
		);
//A34A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A34B65(
		.clk(clk),
			.A(A[34][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1714])
		);
//A35A35
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B35(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[35][BIT_LEN-1:0]),
			.P(mul_result[1715])
		);
//A35A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B36(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1716])
		);
//A35A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B37(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1717])
		);
//A35A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B38(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1718])
		);
//A35A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B39(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1719])
		);
//A35A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B40(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1720])
		);
//A35A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B41(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1721])
		);
//A35A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B42(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1722])
		);
//A35A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B43(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1723])
		);
//A35A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B44(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1724])
		);
//A35A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B45(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1725])
		);
//A35A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B46(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1726])
		);
//A35A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B47(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1727])
		);
//A35A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B48(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1728])
		);
//A35A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B49(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1729])
		);
//A35A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B50(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1730])
		);
//A35A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B51(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1731])
		);
//A35A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B52(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1732])
		);
//A35A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B53(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1733])
		);
//A35A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B54(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1734])
		);
//A35A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B55(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1735])
		);
//A35A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B56(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1736])
		);
//A35A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B57(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1737])
		);
//A35A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B58(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1738])
		);
//A35A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B59(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1739])
		);
//A35A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B60(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1740])
		);
//A35A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B61(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1741])
		);
//A35A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B62(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1742])
		);
//A35A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B63(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1743])
		);
//A35A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B64(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1744])
		);
//A35A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A35B65(
		.clk(clk),
			.A(A[35][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1745])
		);
//A36A36
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B36(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[36][BIT_LEN-1:0]),
			.P(mul_result[1746])
		);
//A36A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B37(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1747])
		);
//A36A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B38(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1748])
		);
//A36A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B39(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1749])
		);
//A36A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B40(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1750])
		);
//A36A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B41(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1751])
		);
//A36A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B42(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1752])
		);
//A36A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B43(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1753])
		);
//A36A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B44(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1754])
		);
//A36A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B45(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1755])
		);
//A36A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B46(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1756])
		);
//A36A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B47(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1757])
		);
//A36A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B48(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1758])
		);
//A36A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B49(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1759])
		);
//A36A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B50(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1760])
		);
//A36A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B51(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1761])
		);
//A36A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B52(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1762])
		);
//A36A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B53(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1763])
		);
//A36A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B54(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1764])
		);
//A36A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B55(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1765])
		);
//A36A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B56(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1766])
		);
//A36A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B57(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1767])
		);
//A36A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B58(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1768])
		);
//A36A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B59(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1769])
		);
//A36A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B60(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1770])
		);
//A36A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B61(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1771])
		);
//A36A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B62(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1772])
		);
//A36A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B63(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1773])
		);
//A36A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B64(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1774])
		);
//A36A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A36B65(
		.clk(clk),
			.A(A[36][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1775])
		);
//A37A37
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B37(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[37][BIT_LEN-1:0]),
			.P(mul_result[1776])
		);
//A37A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B38(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1777])
		);
//A37A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B39(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1778])
		);
//A37A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B40(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1779])
		);
//A37A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B41(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1780])
		);
//A37A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B42(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1781])
		);
//A37A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B43(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1782])
		);
//A37A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B44(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1783])
		);
//A37A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B45(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1784])
		);
//A37A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B46(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1785])
		);
//A37A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B47(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1786])
		);
//A37A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B48(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1787])
		);
//A37A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B49(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1788])
		);
//A37A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B50(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1789])
		);
//A37A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B51(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1790])
		);
//A37A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B52(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1791])
		);
//A37A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B53(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1792])
		);
//A37A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B54(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1793])
		);
//A37A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B55(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1794])
		);
//A37A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B56(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1795])
		);
//A37A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B57(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1796])
		);
//A37A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B58(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1797])
		);
//A37A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B59(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1798])
		);
//A37A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B60(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1799])
		);
//A37A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B61(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1800])
		);
//A37A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B62(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1801])
		);
//A37A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B63(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1802])
		);
//A37A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B64(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1803])
		);
//A37A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A37B65(
		.clk(clk),
			.A(A[37][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1804])
		);
//A38A38
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B38(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[38][BIT_LEN-1:0]),
			.P(mul_result[1805])
		);
//A38A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B39(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1806])
		);
//A38A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B40(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1807])
		);
//A38A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B41(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1808])
		);
//A38A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B42(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1809])
		);
//A38A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B43(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1810])
		);
//A38A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B44(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1811])
		);
//A38A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B45(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1812])
		);
//A38A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B46(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1813])
		);
//A38A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B47(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1814])
		);
//A38A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B48(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1815])
		);
//A38A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B49(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1816])
		);
//A38A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B50(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1817])
		);
//A38A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B51(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1818])
		);
//A38A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B52(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1819])
		);
//A38A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B53(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1820])
		);
//A38A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B54(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1821])
		);
//A38A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B55(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1822])
		);
//A38A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B56(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1823])
		);
//A38A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B57(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1824])
		);
//A38A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B58(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1825])
		);
//A38A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B59(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1826])
		);
//A38A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B60(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1827])
		);
//A38A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B61(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1828])
		);
//A38A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B62(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1829])
		);
//A38A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B63(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1830])
		);
//A38A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B64(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1831])
		);
//A38A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A38B65(
		.clk(clk),
			.A(A[38][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1832])
		);
//A39A39
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B39(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[39][BIT_LEN-1:0]),
			.P(mul_result[1833])
		);
//A39A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B40(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1834])
		);
//A39A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B41(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1835])
		);
//A39A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B42(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1836])
		);
//A39A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B43(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1837])
		);
//A39A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B44(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1838])
		);
//A39A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B45(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1839])
		);
//A39A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B46(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1840])
		);
//A39A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B47(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1841])
		);
//A39A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B48(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1842])
		);
//A39A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B49(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1843])
		);
//A39A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B50(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1844])
		);
//A39A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B51(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1845])
		);
//A39A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B52(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1846])
		);
//A39A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B53(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1847])
		);
//A39A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B54(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1848])
		);
//A39A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B55(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1849])
		);
//A39A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B56(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1850])
		);
//A39A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B57(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1851])
		);
//A39A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B58(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1852])
		);
//A39A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B59(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1853])
		);
//A39A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B60(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1854])
		);
//A39A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B61(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1855])
		);
//A39A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B62(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1856])
		);
//A39A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B63(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1857])
		);
//A39A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B64(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1858])
		);
//A39A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A39B65(
		.clk(clk),
			.A(A[39][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1859])
		);
//A40A40
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B40(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[40][BIT_LEN-1:0]),
			.P(mul_result[1860])
		);
//A40A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B41(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1861])
		);
//A40A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B42(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1862])
		);
//A40A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B43(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1863])
		);
//A40A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B44(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1864])
		);
//A40A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B45(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1865])
		);
//A40A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B46(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1866])
		);
//A40A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B47(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1867])
		);
//A40A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B48(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1868])
		);
//A40A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B49(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1869])
		);
//A40A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B50(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1870])
		);
//A40A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B51(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1871])
		);
//A40A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B52(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1872])
		);
//A40A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B53(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1873])
		);
//A40A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B54(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1874])
		);
//A40A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B55(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1875])
		);
//A40A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B56(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1876])
		);
//A40A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B57(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1877])
		);
//A40A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B58(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1878])
		);
//A40A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B59(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1879])
		);
//A40A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B60(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1880])
		);
//A40A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B61(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1881])
		);
//A40A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B62(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1882])
		);
//A40A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B63(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1883])
		);
//A40A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B64(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1884])
		);
//A40A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A40B65(
		.clk(clk),
			.A(A[40][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1885])
		);
//A41A41
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B41(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[41][BIT_LEN-1:0]),
			.P(mul_result[1886])
		);
//A41A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B42(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1887])
		);
//A41A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B43(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1888])
		);
//A41A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B44(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1889])
		);
//A41A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B45(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1890])
		);
//A41A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B46(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1891])
		);
//A41A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B47(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1892])
		);
//A41A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B48(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1893])
		);
//A41A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B49(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1894])
		);
//A41A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B50(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1895])
		);
//A41A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B51(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1896])
		);
//A41A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B52(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1897])
		);
//A41A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B53(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1898])
		);
//A41A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B54(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1899])
		);
//A41A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B55(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1900])
		);
//A41A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B56(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1901])
		);
//A41A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B57(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1902])
		);
//A41A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B58(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1903])
		);
//A41A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B59(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1904])
		);
//A41A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B60(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1905])
		);
//A41A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B61(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1906])
		);
//A41A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B62(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1907])
		);
//A41A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B63(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1908])
		);
//A41A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B64(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1909])
		);
//A41A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A41B65(
		.clk(clk),
			.A(A[41][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1910])
		);
//A42A42
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B42(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[42][BIT_LEN-1:0]),
			.P(mul_result[1911])
		);
//A42A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B43(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1912])
		);
//A42A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B44(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1913])
		);
//A42A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B45(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1914])
		);
//A42A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B46(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1915])
		);
//A42A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B47(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1916])
		);
//A42A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B48(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1917])
		);
//A42A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B49(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1918])
		);
//A42A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B50(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1919])
		);
//A42A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B51(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1920])
		);
//A42A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B52(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1921])
		);
//A42A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B53(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1922])
		);
//A42A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B54(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1923])
		);
//A42A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B55(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1924])
		);
//A42A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B56(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1925])
		);
//A42A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B57(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1926])
		);
//A42A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B58(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1927])
		);
//A42A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B59(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1928])
		);
//A42A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B60(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1929])
		);
//A42A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B61(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1930])
		);
//A42A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B62(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1931])
		);
//A42A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B63(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1932])
		);
//A42A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B64(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1933])
		);
//A42A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A42B65(
		.clk(clk),
			.A(A[42][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1934])
		);
//A43A43
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B43(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[43][BIT_LEN-1:0]),
			.P(mul_result[1935])
		);
//A43A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B44(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1936])
		);
//A43A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B45(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1937])
		);
//A43A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B46(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1938])
		);
//A43A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B47(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1939])
		);
//A43A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B48(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1940])
		);
//A43A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B49(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1941])
		);
//A43A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B50(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1942])
		);
//A43A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B51(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1943])
		);
//A43A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B52(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1944])
		);
//A43A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B53(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1945])
		);
//A43A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B54(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1946])
		);
//A43A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B55(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1947])
		);
//A43A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B56(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1948])
		);
//A43A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B57(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1949])
		);
//A43A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B58(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1950])
		);
//A43A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B59(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1951])
		);
//A43A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B60(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1952])
		);
//A43A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B61(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1953])
		);
//A43A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B62(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1954])
		);
//A43A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B63(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1955])
		);
//A43A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B64(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1956])
		);
//A43A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A43B65(
		.clk(clk),
			.A(A[43][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1957])
		);
//A44A44
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B44(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[44][BIT_LEN-1:0]),
			.P(mul_result[1958])
		);
//A44A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B45(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1959])
		);
//A44A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B46(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1960])
		);
//A44A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B47(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1961])
		);
//A44A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B48(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1962])
		);
//A44A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B49(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1963])
		);
//A44A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B50(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1964])
		);
//A44A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B51(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1965])
		);
//A44A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B52(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1966])
		);
//A44A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B53(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1967])
		);
//A44A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B54(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1968])
		);
//A44A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B55(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1969])
		);
//A44A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B56(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1970])
		);
//A44A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B57(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1971])
		);
//A44A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B58(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1972])
		);
//A44A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B59(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1973])
		);
//A44A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B60(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1974])
		);
//A44A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B61(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1975])
		);
//A44A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B62(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1976])
		);
//A44A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B63(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1977])
		);
//A44A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B64(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1978])
		);
//A44A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A44B65(
		.clk(clk),
			.A(A[44][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[1979])
		);
//A45A45
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B45(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[45][BIT_LEN-1:0]),
			.P(mul_result[1980])
		);
//A45A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B46(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[1981])
		);
//A45A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B47(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[1982])
		);
//A45A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B48(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[1983])
		);
//A45A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B49(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[1984])
		);
//A45A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B50(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[1985])
		);
//A45A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B51(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[1986])
		);
//A45A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B52(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[1987])
		);
//A45A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B53(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[1988])
		);
//A45A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B54(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[1989])
		);
//A45A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B55(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[1990])
		);
//A45A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B56(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[1991])
		);
//A45A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B57(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[1992])
		);
//A45A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B58(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[1993])
		);
//A45A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B59(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[1994])
		);
//A45A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B60(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[1995])
		);
//A45A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B61(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[1996])
		);
//A45A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B62(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[1997])
		);
//A45A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B63(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[1998])
		);
//A45A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B64(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[1999])
		);
//A45A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A45B65(
		.clk(clk),
			.A(A[45][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2000])
		);
//A46A46
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B46(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[46][BIT_LEN-1:0]),
			.P(mul_result[2001])
		);
//A46A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B47(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[2002])
		);
//A46A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B48(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[2003])
		);
//A46A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B49(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[2004])
		);
//A46A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B50(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[2005])
		);
//A46A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B51(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[2006])
		);
//A46A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B52(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[2007])
		);
//A46A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B53(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2008])
		);
//A46A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B54(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2009])
		);
//A46A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B55(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2010])
		);
//A46A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B56(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2011])
		);
//A46A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B57(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2012])
		);
//A46A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B58(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2013])
		);
//A46A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B59(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2014])
		);
//A46A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B60(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2015])
		);
//A46A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B61(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2016])
		);
//A46A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B62(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2017])
		);
//A46A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B63(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2018])
		);
//A46A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B64(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2019])
		);
//A46A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A46B65(
		.clk(clk),
			.A(A[46][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2020])
		);
//A47A47
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B47(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[47][BIT_LEN-1:0]),
			.P(mul_result[2021])
		);
//A47A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B48(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[2022])
		);
//A47A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B49(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[2023])
		);
//A47A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B50(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[2024])
		);
//A47A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B51(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[2025])
		);
//A47A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B52(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[2026])
		);
//A47A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B53(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2027])
		);
//A47A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B54(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2028])
		);
//A47A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B55(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2029])
		);
//A47A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B56(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2030])
		);
//A47A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B57(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2031])
		);
//A47A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B58(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2032])
		);
//A47A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B59(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2033])
		);
//A47A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B60(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2034])
		);
//A47A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B61(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2035])
		);
//A47A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B62(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2036])
		);
//A47A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B63(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2037])
		);
//A47A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B64(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2038])
		);
//A47A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A47B65(
		.clk(clk),
			.A(A[47][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2039])
		);
//A48A48
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B48(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[48][BIT_LEN-1:0]),
			.P(mul_result[2040])
		);
//A48A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B49(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[2041])
		);
//A48A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B50(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[2042])
		);
//A48A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B51(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[2043])
		);
//A48A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B52(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[2044])
		);
//A48A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B53(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2045])
		);
//A48A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B54(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2046])
		);
//A48A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B55(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2047])
		);
//A48A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B56(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2048])
		);
//A48A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B57(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2049])
		);
//A48A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B58(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2050])
		);
//A48A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B59(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2051])
		);
//A48A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B60(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2052])
		);
//A48A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B61(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2053])
		);
//A48A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B62(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2054])
		);
//A48A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B63(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2055])
		);
//A48A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B64(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2056])
		);
//A48A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A48B65(
		.clk(clk),
			.A(A[48][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2057])
		);
//A49A49
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B49(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[49][BIT_LEN-1:0]),
			.P(mul_result[2058])
		);
//A49A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B50(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[2059])
		);
//A49A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B51(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[2060])
		);
//A49A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B52(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[2061])
		);
//A49A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B53(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2062])
		);
//A49A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B54(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2063])
		);
//A49A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B55(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2064])
		);
//A49A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B56(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2065])
		);
//A49A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B57(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2066])
		);
//A49A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B58(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2067])
		);
//A49A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B59(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2068])
		);
//A49A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B60(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2069])
		);
//A49A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B61(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2070])
		);
//A49A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B62(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2071])
		);
//A49A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B63(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2072])
		);
//A49A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B64(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2073])
		);
//A49A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A49B65(
		.clk(clk),
			.A(A[49][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2074])
		);
//A50A50
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B50(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[50][BIT_LEN-1:0]),
			.P(mul_result[2075])
		);
//A50A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B51(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[2076])
		);
//A50A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B52(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[2077])
		);
//A50A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B53(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2078])
		);
//A50A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B54(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2079])
		);
//A50A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B55(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2080])
		);
//A50A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B56(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2081])
		);
//A50A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B57(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2082])
		);
//A50A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B58(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2083])
		);
//A50A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B59(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2084])
		);
//A50A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B60(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2085])
		);
//A50A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B61(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2086])
		);
//A50A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B62(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2087])
		);
//A50A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B63(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2088])
		);
//A50A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B64(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2089])
		);
//A50A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A50B65(
		.clk(clk),
			.A(A[50][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2090])
		);
//A51A51
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B51(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[51][BIT_LEN-1:0]),
			.P(mul_result[2091])
		);
//A51A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B52(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[2092])
		);
//A51A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B53(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2093])
		);
//A51A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B54(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2094])
		);
//A51A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B55(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2095])
		);
//A51A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B56(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2096])
		);
//A51A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B57(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2097])
		);
//A51A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B58(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2098])
		);
//A51A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B59(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2099])
		);
//A51A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B60(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2100])
		);
//A51A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B61(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2101])
		);
//A51A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B62(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2102])
		);
//A51A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B63(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2103])
		);
//A51A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B64(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2104])
		);
//A51A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A51B65(
		.clk(clk),
			.A(A[51][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2105])
		);
//A52A52
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B52(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[52][BIT_LEN-1:0]),
			.P(mul_result[2106])
		);
//A52A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B53(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2107])
		);
//A52A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B54(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2108])
		);
//A52A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B55(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2109])
		);
//A52A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B56(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2110])
		);
//A52A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B57(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2111])
		);
//A52A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B58(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2112])
		);
//A52A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B59(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2113])
		);
//A52A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B60(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2114])
		);
//A52A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B61(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2115])
		);
//A52A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B62(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2116])
		);
//A52A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B63(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2117])
		);
//A52A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B64(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2118])
		);
//A52A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A52B65(
		.clk(clk),
			.A(A[52][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2119])
		);
//A53A53
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B53(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[53][BIT_LEN-1:0]),
			.P(mul_result[2120])
		);
//A53A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B54(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2121])
		);
//A53A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B55(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2122])
		);
//A53A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B56(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2123])
		);
//A53A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B57(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2124])
		);
//A53A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B58(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2125])
		);
//A53A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B59(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2126])
		);
//A53A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B60(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2127])
		);
//A53A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B61(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2128])
		);
//A53A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B62(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2129])
		);
//A53A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B63(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2130])
		);
//A53A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B64(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2131])
		);
//A53A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A53B65(
		.clk(clk),
			.A(A[53][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2132])
		);
//A54A54
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B54(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[54][BIT_LEN-1:0]),
			.P(mul_result[2133])
		);
//A54A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B55(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2134])
		);
//A54A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B56(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2135])
		);
//A54A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B57(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2136])
		);
//A54A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B58(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2137])
		);
//A54A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B59(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2138])
		);
//A54A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B60(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2139])
		);
//A54A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B61(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2140])
		);
//A54A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B62(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2141])
		);
//A54A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B63(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2142])
		);
//A54A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B64(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2143])
		);
//A54A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A54B65(
		.clk(clk),
			.A(A[54][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2144])
		);
//A55A55
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B55(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[55][BIT_LEN-1:0]),
			.P(mul_result[2145])
		);
//A55A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B56(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2146])
		);
//A55A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B57(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2147])
		);
//A55A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B58(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2148])
		);
//A55A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B59(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2149])
		);
//A55A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B60(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2150])
		);
//A55A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B61(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2151])
		);
//A55A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B62(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2152])
		);
//A55A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B63(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2153])
		);
//A55A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B64(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2154])
		);
//A55A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A55B65(
		.clk(clk),
			.A(A[55][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2155])
		);
//A56A56
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B56(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[56][BIT_LEN-1:0]),
			.P(mul_result[2156])
		);
//A56A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B57(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2157])
		);
//A56A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B58(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2158])
		);
//A56A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B59(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2159])
		);
//A56A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B60(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2160])
		);
//A56A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B61(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2161])
		);
//A56A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B62(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2162])
		);
//A56A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B63(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2163])
		);
//A56A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B64(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2164])
		);
//A56A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A56B65(
		.clk(clk),
			.A(A[56][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2165])
		);
//A57A57
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B57(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[57][BIT_LEN-1:0]),
			.P(mul_result[2166])
		);
//A57A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B58(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2167])
		);
//A57A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B59(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2168])
		);
//A57A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B60(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2169])
		);
//A57A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B61(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2170])
		);
//A57A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B62(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2171])
		);
//A57A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B63(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2172])
		);
//A57A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B64(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2173])
		);
//A57A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A57B65(
		.clk(clk),
			.A(A[57][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2174])
		);
//A58A58
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B58(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[58][BIT_LEN-1:0]),
			.P(mul_result[2175])
		);
//A58A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B59(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2176])
		);
//A58A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B60(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2177])
		);
//A58A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B61(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2178])
		);
//A58A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B62(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2179])
		);
//A58A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B63(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2180])
		);
//A58A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B64(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2181])
		);
//A58A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A58B65(
		.clk(clk),
			.A(A[58][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2182])
		);
//A59A59
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A59B59(
		.clk(clk),
			.A(A[59][BIT_LEN-1:0]),
			.B(B[59][BIT_LEN-1:0]),
			.P(mul_result[2183])
		);
//A59A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A59B60(
		.clk(clk),
			.A(A[59][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2184])
		);
//A59A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A59B61(
		.clk(clk),
			.A(A[59][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2185])
		);
//A59A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A59B62(
		.clk(clk),
			.A(A[59][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2186])
		);
//A59A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A59B63(
		.clk(clk),
			.A(A[59][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2187])
		);
//A59A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A59B64(
		.clk(clk),
			.A(A[59][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2188])
		);
//A59A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A59B65(
		.clk(clk),
			.A(A[59][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2189])
		);
//A60A60
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A60B60(
		.clk(clk),
			.A(A[60][BIT_LEN-1:0]),
			.B(B[60][BIT_LEN-1:0]),
			.P(mul_result[2190])
		);
//A60A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A60B61(
		.clk(clk),
			.A(A[60][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2191])
		);
//A60A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A60B62(
		.clk(clk),
			.A(A[60][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2192])
		);
//A60A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A60B63(
		.clk(clk),
			.A(A[60][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2193])
		);
//A60A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A60B64(
		.clk(clk),
			.A(A[60][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2194])
		);
//A60A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A60B65(
		.clk(clk),
			.A(A[60][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2195])
		);
//A61A61
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A61B61(
		.clk(clk),
			.A(A[61][BIT_LEN-1:0]),
			.B(B[61][BIT_LEN-1:0]),
			.P(mul_result[2196])
		);
//A61A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A61B62(
		.clk(clk),
			.A(A[61][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2197])
		);
//A61A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A61B63(
		.clk(clk),
			.A(A[61][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2198])
		);
//A61A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A61B64(
		.clk(clk),
			.A(A[61][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2199])
		);
//A61A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A61B65(
		.clk(clk),
			.A(A[61][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2200])
		);
//A62A62
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A62B62(
		.clk(clk),
			.A(A[62][BIT_LEN-1:0]),
			.B(B[62][BIT_LEN-1:0]),
			.P(mul_result[2201])
		);
//A62A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A62B63(
		.clk(clk),
			.A(A[62][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2202])
		);
//A62A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A62B64(
		.clk(clk),
			.A(A[62][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2203])
		);
//A62A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A62B65(
		.clk(clk),
			.A(A[62][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2204])
		);
//A63A63
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A63B63(
		.clk(clk),
			.A(A[63][BIT_LEN-1:0]),
			.B(B[63][BIT_LEN-1:0]),
			.P(mul_result[2205])
		);
//A63A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A63B64(
		.clk(clk),
			.A(A[63][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2206])
		);
//A63A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A63B65(
		.clk(clk),
			.A(A[63][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2207])
		);
//A64A64
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A64B64(
		.clk(clk),
			.A(A[64][BIT_LEN-1:0]),
			.B(B[64][BIT_LEN-1:0]),
			.P(mul_result[2208])
		);
//A64A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A64B65(
		.clk(clk),
			.A(A[64][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2209])
		);
//A65A65
multiplier #(.A_BIT_LEN(BIT_LEN),
	.B_BIT_LEN(BIT_LEN)) multiplier_A65B65(
		.clk(clk),
			.A(A[65][BIT_LEN-1:0]),
			.B(B[65][BIT_LEN-1:0]),
			.P(mul_result[2210])
		);
		
		
//MULTIPLIERS register their output therefore we get the results after 1 cycle

// CYCLE 1 starts here
		
		
   //Construct the input wiring thing
   //This is actually the first step of addition (apply the necessary transformations in order to
   //make the addition from x0 + x1 + x1 + x2 + x2 +....+ xn + xn to
   //x0 + 2*x1 + 2*x2 + ... + 2*xn
   //

   //we need to create a grid to facilitate coding + help get it correctly...   
   int ii, jj, index;
      always_comb begin
         for (ii=0; ii<NUM_ELEMENTS*2; ii=ii+1) begin
            for (jj=0; jj<NUM_ELEMENTS*2; jj=jj+1) begin
               grid[ii][jj] = 0;
            end
         end
   	 index = 0;
         for (ii=0; ii<NUM_ELEMENTS; ii=ii+1) begin : grid_row
            for (jj=ii; jj<NUM_ELEMENTS; jj=jj+1) begin : grid_col
               if (jj==ii) begin
               //these are the products that we forward "as is"
               		grid[(ii+jj)][(2*ii)] = {{GRID_PAD_LONG{1'b0}}, mul_result[index][WORD_LEN-1:0]};
               		grid[(ii+jj+1)][((2*ii)+1)] = {{(GRID_PAD_SHORT){1'b0}}, mul_result[index][MUL_OUT_BIT_LEN-1:WORD_LEN]};		
               end
               else begin
               //these are the products that we forward as 2x (ie. left shift by 1)
               		grid[(ii+jj)][(2*ii)] = {{(GRID_PAD_LONG-1){1'b0}}, mul_result[index][WORD_LEN-1:0], 1'b0};
               		grid[(ii+jj+1)][((2*ii)+1)] = {{(GRID_PAD_SHORT-1){1'b0}}, mul_result[index][MUL_OUT_BIT_LEN-1:WORD_LEN], 1'b0};
               end
               index = index +1;
           end
         end
   end
   
   //Calculate all sums (each column of the above constructed grid
   //Remember that the result is in Carry, Sum form (C,S)
   //Remeber #2: the way the grid has been constructed we can use the compressor tree as 
   // provided, however bear in mind that now the maximum number of values to be added is not
   // (2*NUM_ELEMENTS)-1 but NUM_ELEMENTS
       
   genvar i;
   generate
      // The first and last columns have only one entry, return in S
      always_ff @(posedge clk) begin
         Cout[0][OUT_BIT_LEN-1:0]                  <= '0;
         Cout[(NUM_ELEMENTS*2)-1][OUT_BIT_LEN-1:0] <= '0;

         S[0][OUT_BIT_LEN-1:0] <= grid[0][0][OUT_BIT_LEN-1:0];

         S[(NUM_ELEMENTS*2)-1][OUT_BIT_LEN-1:0] <= grid[(NUM_ELEMENTS*2)-1][(NUM_ELEMENTS*2)-1][OUT_BIT_LEN-1:0];
      end

      // Loop through grid parallelogram
      // The number of elements increases up to the midpoint then decreases
      // Starting grid row is 0 for the first half, decreases by 2 thereafter
      // Instantiate compressor tree per column
      for (i=1; i<(NUM_ELEMENTS*2)-1; i=i+1) begin : col_sums
         localparam integer CUR_ELEMENTS = (i < NUM_ELEMENTS) ? (i+1) : ((NUM_ELEMENTS*2) - i);
         localparam integer GRID_INDEX   = (i < NUM_ELEMENTS) ? 0 : (((i - NUM_ELEMENTS) * 2) + 1);

         logic [OUT_BIT_LEN-1:0] Cout_col;
         logic [OUT_BIT_LEN-1:0] S_col; 

         compressor_tree_3_to_2 #(.NUM_ELEMENTS(CUR_ELEMENTS),
                                  .BIT_LEN(OUT_BIT_LEN)
                                 )
            compressor_tree_3_to_2 (
               .terms(grid[i][GRID_INDEX:(GRID_INDEX + CUR_ELEMENTS - 1)]),
               .C(Cout_col),
               .S(S_col)
            );

         always_ff @(posedge clk) begin
            Cout[i][OUT_BIT_LEN-1:0] <= Cout_col[OUT_BIT_LEN-1:0];
            S[i][OUT_BIT_LEN-1:0]    <= S_col[OUT_BIT_LEN-1:0];
         end
      end
   endgenerate   

//CYCLE 2 

// We get the results from the adder trees in C,S form and make the final 
//carry propagate addition
   
	// Carry propogate add each column in grid
	// Partially reduce adding neighbor carries
	always_comb begin
		for (int k = 0; k < NUM_ELEMENTS*2; k = k+1) begin
			//CPA each Cout and S of the CSA to get final result
			//remember each Cout and S are OUT_BIT_LEN bits long and therefore each grid sum is OUT_BIT_LEN+1 bits long
			grid_sum[k] = Cout[k] + S[k];
		end

		//In the reduced_grid_sum all numbers are BIT_LEN (17) bits long
		reduced_grid_sum[0] = {{(BIT_LEN-WORD_LEN){1'b0}}, grid_sum[0][WORD_LEN-1:0]};

		for (int k=1; k<(NUM_ELEMENTS*2)-1; k=k+1) begin
			//Consider each coefficient is BIT_LEN bits long.
			//Add the carry from the previous coefficient.
			reduced_grid_sum[k] = {{(BIT_LEN-WORD_LEN){1'b0}}, grid_sum[k][WORD_LEN-1:0]} + {{(BIT_LEN-(OUT_BIT_LEN-WORD_LEN))-1{1'b0}}, grid_sum[k-1][OUT_BIT_LEN:WORD_LEN]};
		end
		reduced_grid_sum[(NUM_ELEMENTS*2)-1] = grid_sum[(NUM_ELEMENTS*2)-1][BIT_LEN-1:0] +  {{(BIT_LEN-(OUT_BIT_LEN-WORD_LEN))-1{1'b0}}, grid_sum[(NUM_ELEMENTS*2)-2][OUT_BIT_LEN:WORD_LEN]};
	end
	
	//register outputs
	always_ff @(posedge clk) begin
   		for (int k = 0; k < NUM_ELEMENTS*2; k = k+1) begin
   			reduced_output[k] <= reduced_grid_sum[k];
   		end
 	end
	
	
	
	
endmodule
   

